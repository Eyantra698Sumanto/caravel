magic
tech sky130A
magscale 1 2
timestamp 1685569056
<< checkpaint >>
rect -194 868 20158 18716
<< viali >>
rect 1593 17289 1627 17323
rect 4169 17289 4203 17323
rect 5089 17289 5123 17323
rect 6929 17289 6963 17323
rect 15761 17289 15795 17323
rect 18061 17289 18095 17323
rect 4629 17221 4663 17255
rect 12449 17221 12483 17255
rect 1501 17153 1535 17187
rect 2145 17153 2179 17187
rect 4077 17153 4111 17187
rect 4537 17153 4571 17187
rect 4997 17153 5031 17187
rect 5181 17153 5215 17187
rect 6653 17153 6687 17187
rect 9781 17153 9815 17187
rect 10149 17153 10183 17187
rect 15669 17153 15703 17187
rect 17785 17153 17819 17187
rect 5365 17085 5399 17119
rect 1961 17017 1995 17051
rect 4813 17017 4847 17051
rect 12633 17017 12667 17051
rect 9965 16949 9999 16983
rect 10241 16949 10275 16983
rect 4445 16745 4479 16779
rect 14473 16745 14507 16779
rect 16957 16745 16991 16779
rect 18245 16745 18279 16779
rect 17141 16677 17175 16711
rect 14105 16609 14139 16643
rect 4169 16541 4203 16575
rect 10057 16541 10091 16575
rect 12817 16541 12851 16575
rect 14289 16541 14323 16575
rect 16773 16473 16807 16507
rect 18153 16473 18187 16507
rect 4629 16405 4663 16439
rect 10149 16405 10183 16439
rect 12909 16405 12943 16439
rect 16973 16405 17007 16439
rect 3249 16201 3283 16235
rect 12909 16201 12943 16235
rect 14933 16201 14967 16235
rect 13461 16133 13495 16167
rect 3157 16065 3191 16099
rect 3341 16065 3375 16099
rect 7481 16065 7515 16099
rect 7665 16065 7699 16099
rect 15025 16065 15059 16099
rect 15209 16065 15243 16099
rect 15485 16065 15519 16099
rect 15761 16065 15795 16099
rect 16865 16065 16899 16099
rect 18245 16065 18279 16099
rect 7757 15997 7791 16031
rect 8033 15997 8067 16031
rect 12633 15997 12667 16031
rect 12725 15997 12759 16031
rect 13001 15997 13035 16031
rect 13093 15997 13127 16031
rect 13185 15997 13219 16031
rect 16957 15997 16991 16031
rect 2973 15929 3007 15963
rect 3525 15861 3559 15895
rect 7481 15861 7515 15895
rect 9505 15861 9539 15895
rect 12449 15861 12483 15895
rect 15025 15861 15059 15895
rect 15577 15861 15611 15895
rect 15853 15861 15887 15895
rect 17233 15861 17267 15895
rect 18429 15861 18463 15895
rect 4997 15657 5031 15691
rect 13461 15657 13495 15691
rect 12449 15589 12483 15623
rect 4537 15521 4571 15555
rect 10701 15521 10735 15555
rect 15853 15521 15887 15555
rect 1501 15453 1535 15487
rect 13645 15453 13679 15487
rect 13921 15453 13955 15487
rect 14105 15453 14139 15487
rect 3801 15385 3835 15419
rect 4813 15385 4847 15419
rect 10977 15385 11011 15419
rect 14381 15385 14415 15419
rect 1593 15317 1627 15351
rect 5013 15317 5047 15351
rect 5181 15317 5215 15351
rect 13829 15317 13863 15351
rect 11805 15113 11839 15147
rect 11897 15113 11931 15147
rect 11989 15113 12023 15147
rect 15117 15045 15151 15079
rect 11161 14977 11195 15011
rect 11253 14977 11287 15011
rect 12357 14977 12391 15011
rect 14749 14977 14783 15011
rect 15209 14977 15243 15011
rect 17693 14977 17727 15011
rect 17877 14977 17911 15011
rect 11621 14909 11655 14943
rect 12633 14909 12667 14943
rect 12173 14841 12207 14875
rect 17325 14841 17359 14875
rect 14105 14773 14139 14807
rect 15301 14773 15335 14807
rect 17693 14773 17727 14807
rect 6561 14569 6595 14603
rect 12265 14569 12299 14603
rect 17049 14501 17083 14535
rect 6285 14433 6319 14467
rect 11897 14433 11931 14467
rect 17141 14433 17175 14467
rect 3157 14365 3191 14399
rect 6193 14365 6227 14399
rect 6469 14365 6503 14399
rect 11805 14365 11839 14399
rect 13645 14365 13679 14399
rect 17049 14365 17083 14399
rect 2789 14297 2823 14331
rect 12081 14297 12115 14331
rect 17325 14297 17359 14331
rect 2973 14229 3007 14263
rect 3065 14229 3099 14263
rect 3341 14229 3375 14263
rect 12281 14229 12315 14263
rect 12449 14229 12483 14263
rect 13461 14229 13495 14263
rect 2513 13889 2547 13923
rect 4445 13889 4479 13923
rect 6837 13889 6871 13923
rect 2237 13821 2271 13855
rect 2789 13821 2823 13855
rect 4261 13821 4295 13855
rect 4537 13821 4571 13855
rect 7205 13821 7239 13855
rect 7481 13821 7515 13855
rect 8953 13821 8987 13855
rect 13829 13821 13863 13855
rect 15577 13821 15611 13855
rect 7021 13685 7055 13719
rect 14092 13685 14126 13719
rect 17325 13481 17359 13515
rect 15301 13413 15335 13447
rect 15853 13345 15887 13379
rect 2145 13277 2179 13311
rect 2421 13277 2455 13311
rect 2605 13277 2639 13311
rect 2973 13277 3007 13311
rect 3157 13277 3191 13311
rect 3801 13277 3835 13311
rect 6285 13277 6319 13311
rect 10609 13277 10643 13311
rect 13737 13277 13771 13311
rect 14473 13277 14507 13311
rect 15117 13277 15151 13311
rect 15577 13277 15611 13311
rect 2329 13209 2363 13243
rect 13829 13209 13863 13243
rect 14105 13209 14139 13243
rect 3893 13141 3927 13175
rect 6377 13141 6411 13175
rect 10701 13141 10735 13175
rect 14289 13141 14323 13175
rect 14381 13141 14415 13175
rect 14657 13141 14691 13175
rect 1409 12937 1443 12971
rect 18245 12937 18279 12971
rect 1593 12801 1627 12835
rect 7205 12801 7239 12835
rect 7665 12801 7699 12835
rect 18153 12801 18187 12835
rect 2605 12733 2639 12767
rect 2881 12733 2915 12767
rect 7297 12733 7331 12767
rect 7941 12733 7975 12767
rect 9413 12733 9447 12767
rect 14749 12733 14783 12767
rect 15025 12733 15059 12767
rect 4353 12597 4387 12631
rect 7573 12597 7607 12631
rect 16497 12597 16531 12631
rect 2053 12393 2087 12427
rect 8953 12393 8987 12427
rect 9965 12393 9999 12427
rect 10701 12393 10735 12427
rect 14473 12393 14507 12427
rect 2973 12325 3007 12359
rect 10885 12325 10919 12359
rect 3249 12257 3283 12291
rect 6285 12257 6319 12291
rect 6377 12257 6411 12291
rect 6561 12257 6595 12291
rect 9229 12257 9263 12291
rect 9413 12257 9447 12291
rect 9597 12257 9631 12291
rect 2237 12189 2271 12223
rect 2513 12189 2547 12223
rect 3157 12189 3191 12223
rect 3341 12189 3375 12223
rect 3433 12189 3467 12223
rect 6469 12189 6503 12223
rect 7297 12189 7331 12223
rect 9137 12189 9171 12223
rect 9321 12189 9355 12223
rect 9781 12189 9815 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 10333 12121 10367 12155
rect 2421 12053 2455 12087
rect 6101 12053 6135 12087
rect 7389 12053 7423 12087
rect 10710 12053 10744 12087
rect 6377 11849 6411 11883
rect 14013 11849 14047 11883
rect 1961 11713 1995 11747
rect 2145 11713 2179 11747
rect 2329 11713 2363 11747
rect 2605 11713 2639 11747
rect 2798 11713 2832 11747
rect 6653 11713 6687 11747
rect 7021 11713 7055 11747
rect 10421 11713 10455 11747
rect 14197 11713 14231 11747
rect 3433 11645 3467 11679
rect 6561 11645 6595 11679
rect 6745 11645 6779 11679
rect 6837 11645 6871 11679
rect 10517 11645 10551 11679
rect 10609 11645 10643 11679
rect 10701 11645 10735 11679
rect 12265 11645 12299 11679
rect 7481 11577 7515 11611
rect 7113 11509 7147 11543
rect 10241 11509 10275 11543
rect 12528 11509 12562 11543
rect 14381 11509 14415 11543
rect 3801 11305 3835 11339
rect 4537 11305 4571 11339
rect 8953 11305 8987 11339
rect 18521 11305 18555 11339
rect 9965 11237 9999 11271
rect 10057 11237 10091 11271
rect 15853 11237 15887 11271
rect 4077 11169 4111 11203
rect 4445 11169 4479 11203
rect 4813 11169 4847 11203
rect 4905 11169 4939 11203
rect 9229 11169 9263 11203
rect 14381 11169 14415 11203
rect 18153 11169 18187 11203
rect 3985 11101 4019 11135
rect 4721 11101 4755 11135
rect 4997 11101 5031 11135
rect 9137 11101 9171 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 10333 11101 10367 11135
rect 14105 11101 14139 11135
rect 18337 11101 18371 11135
rect 9597 11033 9631 11067
rect 10609 11033 10643 11067
rect 12357 11033 12391 11067
rect 4261 10965 4295 10999
rect 4353 10965 4387 10999
rect 7573 10761 7607 10795
rect 2789 10693 2823 10727
rect 17233 10693 17267 10727
rect 17417 10693 17451 10727
rect 17969 10693 18003 10727
rect 18185 10693 18219 10727
rect 2697 10625 2731 10659
rect 3617 10625 3651 10659
rect 7481 10625 7515 10659
rect 17693 10625 17727 10659
rect 14933 10557 14967 10591
rect 15209 10489 15243 10523
rect 3709 10421 3743 10455
rect 15393 10421 15427 10455
rect 17417 10421 17451 10455
rect 18153 10421 18187 10455
rect 18337 10421 18371 10455
rect 15669 10217 15703 10251
rect 17049 10149 17083 10183
rect 4537 10081 4571 10115
rect 4629 10081 4663 10115
rect 4813 10081 4847 10115
rect 7389 10081 7423 10115
rect 7481 10081 7515 10115
rect 7665 10081 7699 10115
rect 10609 10081 10643 10115
rect 16037 10081 16071 10115
rect 4721 10013 4755 10047
rect 4997 10013 5031 10047
rect 7573 10013 7607 10047
rect 15853 10013 15887 10047
rect 15945 10013 15979 10047
rect 16129 10013 16163 10047
rect 17325 10013 17359 10047
rect 17417 10013 17451 10047
rect 5273 9945 5307 9979
rect 10885 9945 10919 9979
rect 18153 9945 18187 9979
rect 4353 9877 4387 9911
rect 6745 9877 6779 9911
rect 7205 9877 7239 9911
rect 12357 9877 12391 9911
rect 17233 9877 17267 9911
rect 17601 9877 17635 9911
rect 18245 9877 18279 9911
rect 1777 9605 1811 9639
rect 14289 9605 14323 9639
rect 14473 9605 14507 9639
rect 1685 9537 1719 9571
rect 5181 9537 5215 9571
rect 8585 9537 8619 9571
rect 12265 9537 12299 9571
rect 13461 9537 13495 9571
rect 14565 9537 14599 9571
rect 6469 9469 6503 9503
rect 6745 9469 6779 9503
rect 8217 9469 8251 9503
rect 8861 9469 8895 9503
rect 14289 9401 14323 9435
rect 5273 9333 5307 9367
rect 10333 9333 10367 9367
rect 12357 9333 12391 9367
rect 13645 9333 13679 9367
rect 13921 9129 13955 9163
rect 6929 9061 6963 9095
rect 7665 9061 7699 9095
rect 6770 8993 6804 9027
rect 8125 8993 8159 9027
rect 8217 8993 8251 9027
rect 1501 8925 1535 8959
rect 6285 8925 6319 8959
rect 6653 8925 6687 8959
rect 8953 8925 8987 8959
rect 9229 8925 9263 8959
rect 12173 8925 12207 8959
rect 14933 8925 14967 8959
rect 8033 8857 8067 8891
rect 9321 8857 9355 8891
rect 12449 8857 12483 8891
rect 15761 8857 15795 8891
rect 1593 8789 1627 8823
rect 6561 8789 6595 8823
rect 9137 8789 9171 8823
rect 9505 8789 9539 8823
rect 3801 8585 3835 8619
rect 10609 8585 10643 8619
rect 13737 8585 13771 8619
rect 3433 8449 3467 8483
rect 3617 8449 3651 8483
rect 6377 8449 6411 8483
rect 7297 8449 7331 8483
rect 10517 8449 10551 8483
rect 17693 8449 17727 8483
rect 6561 8381 6595 8415
rect 7021 8381 7055 8415
rect 7414 8381 7448 8415
rect 7573 8381 7607 8415
rect 13921 8381 13955 8415
rect 14013 8381 14047 8415
rect 14105 8381 14139 8415
rect 14197 8381 14231 8415
rect 8217 8313 8251 8347
rect 17969 8313 18003 8347
rect 18153 8313 18187 8347
rect 6285 8041 6319 8075
rect 11069 8041 11103 8075
rect 2881 7973 2915 8007
rect 10149 7973 10183 8007
rect 10241 7905 10275 7939
rect 2789 7837 2823 7871
rect 6469 7837 6503 7871
rect 6745 7837 6779 7871
rect 10977 7837 11011 7871
rect 9781 7769 9815 7803
rect 6653 7701 6687 7735
rect 11989 7497 12023 7531
rect 5457 7361 5491 7395
rect 5917 7361 5951 7395
rect 6101 7361 6135 7395
rect 6193 7361 6227 7395
rect 6837 7361 6871 7395
rect 7665 7361 7699 7395
rect 12173 7361 12207 7395
rect 12449 7361 12483 7395
rect 17877 7361 17911 7395
rect 5549 7293 5583 7327
rect 6561 7293 6595 7327
rect 6653 7293 6687 7327
rect 6745 7293 6779 7327
rect 12357 7293 12391 7327
rect 5825 7225 5859 7259
rect 5917 7157 5951 7191
rect 6377 7157 6411 7191
rect 7849 7157 7883 7191
rect 17969 7157 18003 7191
rect 17417 6817 17451 6851
rect 17325 6749 17359 6783
rect 17969 6749 18003 6783
rect 18061 6681 18095 6715
rect 6193 6409 6227 6443
rect 14013 6409 14047 6443
rect 3433 6341 3467 6375
rect 4721 6341 4755 6375
rect 1501 6273 1535 6307
rect 1961 6273 1995 6307
rect 2513 6273 2547 6307
rect 2789 6273 2823 6307
rect 2973 6273 3007 6307
rect 3249 6273 3283 6307
rect 3525 6273 3559 6307
rect 3985 6273 4019 6307
rect 4445 6273 4479 6307
rect 6561 6273 6595 6307
rect 7573 6273 7607 6307
rect 13737 6273 13771 6307
rect 18245 6273 18279 6307
rect 2329 6205 2363 6239
rect 6653 6205 6687 6239
rect 7849 6205 7883 6239
rect 14013 6205 14047 6239
rect 2053 6137 2087 6171
rect 3065 6137 3099 6171
rect 18429 6137 18463 6171
rect 1593 6069 1627 6103
rect 4169 6069 4203 6103
rect 6929 6069 6963 6103
rect 9321 6069 9355 6103
rect 13829 6069 13863 6103
rect 3985 5865 4019 5899
rect 7389 5865 7423 5899
rect 10149 5865 10183 5899
rect 15669 5865 15703 5899
rect 8033 5797 8067 5831
rect 5733 5729 5767 5763
rect 7573 5729 7607 5763
rect 9689 5729 9723 5763
rect 11989 5729 12023 5763
rect 12081 5729 12115 5763
rect 3985 5661 4019 5695
rect 4169 5661 4203 5695
rect 5457 5661 5491 5695
rect 7665 5661 7699 5695
rect 7757 5661 7791 5695
rect 7849 5661 7883 5695
rect 9781 5661 9815 5695
rect 12173 5661 12207 5695
rect 12265 5661 12299 5695
rect 15485 5661 15519 5695
rect 8217 5593 8251 5627
rect 8585 5593 8619 5627
rect 7205 5525 7239 5559
rect 8309 5525 8343 5559
rect 8401 5525 8435 5559
rect 11805 5525 11839 5559
rect 1869 5321 1903 5355
rect 11713 5321 11747 5355
rect 15853 5321 15887 5355
rect 1777 5253 1811 5287
rect 3985 5253 4019 5287
rect 7665 5253 7699 5287
rect 7849 5253 7883 5287
rect 12265 5253 12299 5287
rect 15761 5253 15795 5287
rect 2421 5185 2455 5219
rect 3709 5185 3743 5219
rect 7481 5185 7515 5219
rect 7573 5185 7607 5219
rect 11805 5185 11839 5219
rect 11897 5185 11931 5219
rect 12173 5185 12207 5219
rect 16037 5185 16071 5219
rect 2053 5117 2087 5151
rect 2513 5117 2547 5151
rect 5457 5117 5491 5151
rect 7297 5049 7331 5083
rect 11529 5049 11563 5083
rect 16221 5049 16255 5083
rect 1409 4981 1443 5015
rect 2789 4981 2823 5015
rect 12081 4981 12115 5015
rect 3157 4777 3191 4811
rect 5273 4777 5307 4811
rect 7389 4777 7423 4811
rect 9597 4777 9631 4811
rect 16957 4777 16991 4811
rect 1409 4641 1443 4675
rect 1685 4641 1719 4675
rect 10057 4641 10091 4675
rect 11897 4641 11931 4675
rect 15485 4641 15519 4675
rect 4261 4573 4295 4607
rect 6009 4573 6043 4607
rect 6745 4573 6779 4607
rect 7021 4573 7055 4607
rect 9781 4573 9815 4607
rect 9873 4573 9907 4607
rect 9966 4573 10000 4607
rect 11621 4573 11655 4607
rect 15209 4573 15243 4607
rect 3985 4505 4019 4539
rect 4353 4505 4387 4539
rect 4721 4505 4755 4539
rect 5089 4437 5123 4471
rect 7389 4437 7423 4471
rect 7573 4437 7607 4471
rect 13369 4437 13403 4471
rect 2355 4233 2389 4267
rect 5825 4233 5859 4267
rect 18245 4233 18279 4267
rect 18429 4233 18463 4267
rect 2145 4165 2179 4199
rect 18061 4165 18095 4199
rect 1501 4097 1535 4131
rect 1685 4097 1719 4131
rect 1961 4097 1995 4131
rect 4077 4097 4111 4131
rect 7573 4097 7607 4131
rect 8217 4097 8251 4131
rect 16681 4097 16715 4131
rect 1777 4029 1811 4063
rect 4353 4029 4387 4063
rect 8309 4029 8343 4063
rect 11529 4029 11563 4063
rect 11805 4029 11839 4063
rect 1869 3961 1903 3995
rect 2513 3961 2547 3995
rect 8585 3961 8619 3995
rect 16957 3961 16991 3995
rect 17417 3961 17451 3995
rect 2329 3893 2363 3927
rect 7389 3893 7423 3927
rect 13277 3893 13311 3927
rect 17141 3893 17175 3927
rect 18245 3893 18279 3927
rect 1593 3689 1627 3723
rect 4629 3689 4663 3723
rect 14822 3689 14856 3723
rect 17509 3689 17543 3723
rect 18245 3689 18279 3723
rect 1501 3621 1535 3655
rect 3893 3621 3927 3655
rect 5825 3621 5859 3655
rect 11161 3621 11195 3655
rect 14933 3621 14967 3655
rect 1685 3553 1719 3587
rect 4445 3553 4479 3587
rect 5457 3553 5491 3587
rect 10977 3553 11011 3587
rect 11805 3553 11839 3587
rect 15025 3553 15059 3587
rect 15117 3553 15151 3587
rect 15485 3553 15519 3587
rect 1409 3485 1443 3519
rect 1777 3485 1811 3519
rect 8953 3485 8987 3519
rect 11069 3485 11103 3519
rect 11897 3485 11931 3519
rect 12265 3485 12299 3519
rect 12541 3485 12575 3519
rect 14657 3485 14691 3519
rect 17417 3485 17451 3519
rect 3893 3417 3927 3451
rect 4353 3417 4387 3451
rect 9229 3417 9263 3451
rect 15761 3417 15795 3451
rect 18153 3417 18187 3451
rect 1869 3349 1903 3383
rect 5917 3349 5951 3383
rect 17233 3349 17267 3383
rect 6577 3145 6611 3179
rect 6745 3145 6779 3179
rect 9689 3145 9723 3179
rect 10517 3145 10551 3179
rect 13185 3145 13219 3179
rect 16329 3145 16363 3179
rect 16497 3145 16531 3179
rect 1501 3077 1535 3111
rect 6377 3077 6411 3111
rect 16129 3077 16163 3111
rect 9505 3009 9539 3043
rect 10701 3009 10735 3043
rect 10977 3009 11011 3043
rect 11713 3009 11747 3043
rect 13093 3009 13127 3043
rect 14841 3009 14875 3043
rect 15301 3009 15335 3043
rect 17141 3009 17175 3043
rect 17417 3009 17451 3043
rect 11621 2941 11655 2975
rect 16957 2941 16991 2975
rect 17233 2941 17267 2975
rect 17325 2941 17359 2975
rect 12081 2873 12115 2907
rect 15485 2873 15519 2907
rect 1593 2805 1627 2839
rect 6561 2805 6595 2839
rect 10885 2805 10919 2839
rect 15117 2805 15151 2839
rect 16313 2805 16347 2839
rect 6101 2601 6135 2635
rect 11897 2601 11931 2635
rect 18337 2601 18371 2635
rect 9137 2533 9171 2567
rect 9321 2465 9355 2499
rect 1501 2397 1535 2431
rect 5917 2397 5951 2431
rect 8401 2397 8435 2431
rect 9045 2397 9079 2431
rect 11345 2397 11379 2431
rect 11713 2397 11747 2431
rect 14381 2397 14415 2431
rect 17601 2397 17635 2431
rect 18521 2397 18555 2431
rect 2789 2329 2823 2363
rect 9597 2329 9631 2363
rect 1593 2261 1627 2295
rect 2881 2261 2915 2295
rect 8493 2261 8527 2295
rect 14473 2261 14507 2295
rect 17693 2261 17727 2295
<< metal1 >>
rect 1104 17434 18860 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 7610 17434
rect 7662 17382 7674 17434
rect 7726 17382 7738 17434
rect 7790 17382 7802 17434
rect 7854 17382 7866 17434
rect 7918 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 17610 17434
rect 17662 17382 17674 17434
rect 17726 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 18860 17434
rect 1104 17360 18860 17382
rect 1578 17280 1584 17332
rect 1636 17280 1642 17332
rect 4154 17280 4160 17332
rect 4212 17280 4218 17332
rect 5077 17323 5135 17329
rect 5077 17320 5089 17323
rect 4540 17292 5089 17320
rect 658 17212 664 17264
rect 716 17252 722 17264
rect 716 17224 2176 17252
rect 716 17212 722 17224
rect 1486 17144 1492 17196
rect 1544 17144 1550 17196
rect 2148 17193 2176 17224
rect 3050 17212 3056 17264
rect 3108 17252 3114 17264
rect 4540 17252 4568 17292
rect 5077 17289 5089 17292
rect 5123 17289 5135 17323
rect 5077 17283 5135 17289
rect 6454 17280 6460 17332
rect 6512 17320 6518 17332
rect 6917 17323 6975 17329
rect 6917 17320 6929 17323
rect 6512 17292 6929 17320
rect 6512 17280 6518 17292
rect 6917 17289 6929 17292
rect 6963 17289 6975 17323
rect 10870 17320 10876 17332
rect 6917 17283 6975 17289
rect 8496 17292 10876 17320
rect 3108 17224 4568 17252
rect 4617 17255 4675 17261
rect 3108 17212 3114 17224
rect 4617 17221 4629 17255
rect 4663 17252 4675 17255
rect 8496 17252 8524 17292
rect 10870 17280 10876 17292
rect 10928 17280 10934 17332
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 15749 17323 15807 17329
rect 15749 17320 15761 17323
rect 15528 17292 15761 17320
rect 15528 17280 15534 17292
rect 15749 17289 15761 17292
rect 15795 17289 15807 17323
rect 15749 17283 15807 17289
rect 17954 17280 17960 17332
rect 18012 17320 18018 17332
rect 18049 17323 18107 17329
rect 18049 17320 18061 17323
rect 18012 17292 18061 17320
rect 18012 17280 18018 17292
rect 18049 17289 18061 17292
rect 18095 17289 18107 17323
rect 18049 17283 18107 17289
rect 4663 17224 8524 17252
rect 8588 17224 10180 17252
rect 4663 17221 4675 17224
rect 4617 17215 4675 17221
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17153 2191 17187
rect 2133 17147 2191 17153
rect 4062 17144 4068 17196
rect 4120 17144 4126 17196
rect 4522 17144 4528 17196
rect 4580 17144 4586 17196
rect 4985 17187 5043 17193
rect 4985 17184 4997 17187
rect 4724 17156 4997 17184
rect 1949 17051 2007 17057
rect 1949 17017 1961 17051
rect 1995 17017 2007 17051
rect 1949 17011 2007 17017
rect 1964 16980 1992 17011
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 4724 17048 4752 17156
rect 4985 17153 4997 17156
rect 5031 17153 5043 17187
rect 4985 17147 5043 17153
rect 5169 17187 5227 17193
rect 5169 17153 5181 17187
rect 5215 17184 5227 17187
rect 6270 17184 6276 17196
rect 5215 17156 6276 17184
rect 5215 17153 5227 17156
rect 5169 17147 5227 17153
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 6638 17144 6644 17196
rect 6696 17144 6702 17196
rect 8588 17184 8616 17224
rect 7392 17156 8616 17184
rect 5350 17076 5356 17128
rect 5408 17076 5414 17128
rect 3016 17020 4752 17048
rect 4801 17051 4859 17057
rect 3016 17008 3022 17020
rect 4801 17017 4813 17051
rect 4847 17048 4859 17051
rect 6454 17048 6460 17060
rect 4847 17020 6460 17048
rect 4847 17017 4859 17020
rect 4801 17011 4859 17017
rect 6454 17008 6460 17020
rect 6512 17008 6518 17060
rect 4338 16980 4344 16992
rect 1964 16952 4344 16980
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 4522 16940 4528 16992
rect 4580 16980 4586 16992
rect 7392 16980 7420 17156
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 10152 17193 10180 17224
rect 12250 17212 12256 17264
rect 12308 17252 12314 17264
rect 12437 17255 12495 17261
rect 12437 17252 12449 17255
rect 12308 17224 12449 17252
rect 12308 17212 12314 17224
rect 12437 17221 12449 17224
rect 12483 17221 12495 17255
rect 12437 17215 12495 17221
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 9732 17156 9781 17184
rect 9732 17144 9738 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 13998 17184 14004 17196
rect 10183 17156 14004 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 15657 17187 15715 17193
rect 15657 17153 15669 17187
rect 15703 17184 15715 17187
rect 15930 17184 15936 17196
rect 15703 17156 15936 17184
rect 15703 17153 15715 17156
rect 15657 17147 15715 17153
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 16724 17156 17785 17184
rect 16724 17144 16730 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 17773 17147 17831 17153
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 14918 17116 14924 17128
rect 8352 17088 14924 17116
rect 8352 17076 8358 17088
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 12621 17051 12679 17057
rect 12621 17017 12633 17051
rect 12667 17048 12679 17051
rect 15194 17048 15200 17060
rect 12667 17020 15200 17048
rect 12667 17017 12679 17020
rect 12621 17011 12679 17017
rect 15194 17008 15200 17020
rect 15252 17008 15258 17060
rect 4580 16952 7420 16980
rect 4580 16940 4586 16952
rect 9950 16940 9956 16992
rect 10008 16940 10014 16992
rect 10229 16983 10287 16989
rect 10229 16949 10241 16983
rect 10275 16980 10287 16983
rect 10410 16980 10416 16992
rect 10275 16952 10416 16980
rect 10275 16949 10287 16952
rect 10229 16943 10287 16949
rect 10410 16940 10416 16952
rect 10468 16940 10474 16992
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 13538 16980 13544 16992
rect 12860 16952 13544 16980
rect 12860 16940 12866 16952
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 1104 16890 18860 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 6950 16890
rect 7002 16838 7014 16890
rect 7066 16838 7078 16890
rect 7130 16838 7142 16890
rect 7194 16838 7206 16890
rect 7258 16838 11950 16890
rect 12002 16838 12014 16890
rect 12066 16838 12078 16890
rect 12130 16838 12142 16890
rect 12194 16838 12206 16890
rect 12258 16838 16950 16890
rect 17002 16838 17014 16890
rect 17066 16838 17078 16890
rect 17130 16838 17142 16890
rect 17194 16838 17206 16890
rect 17258 16838 18860 16890
rect 1104 16816 18860 16838
rect 4433 16779 4491 16785
rect 4433 16745 4445 16779
rect 4479 16776 4491 16779
rect 9214 16776 9220 16788
rect 4479 16748 9220 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 9214 16736 9220 16748
rect 9272 16736 9278 16788
rect 9306 16736 9312 16788
rect 9364 16776 9370 16788
rect 14461 16779 14519 16785
rect 14461 16776 14473 16779
rect 9364 16748 14473 16776
rect 9364 16736 9370 16748
rect 14461 16745 14473 16748
rect 14507 16745 14519 16779
rect 14461 16739 14519 16745
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16945 16779 17003 16785
rect 16945 16776 16957 16779
rect 16356 16748 16957 16776
rect 16356 16736 16362 16748
rect 16945 16745 16957 16748
rect 16991 16745 17003 16779
rect 16945 16739 17003 16745
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 18233 16779 18291 16785
rect 18233 16776 18245 16779
rect 18104 16748 18245 16776
rect 18104 16736 18110 16748
rect 18233 16745 18245 16748
rect 18279 16745 18291 16779
rect 18233 16739 18291 16745
rect 4338 16668 4344 16720
rect 4396 16708 4402 16720
rect 6914 16708 6920 16720
rect 4396 16680 6920 16708
rect 4396 16668 4402 16680
rect 6914 16668 6920 16680
rect 6972 16668 6978 16720
rect 17129 16711 17187 16717
rect 17129 16677 17141 16711
rect 17175 16708 17187 16711
rect 17954 16708 17960 16720
rect 17175 16680 17960 16708
rect 17175 16677 17187 16680
rect 17129 16671 17187 16677
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 8294 16640 8300 16652
rect 4172 16612 8300 16640
rect 4172 16581 4200 16612
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 11790 16600 11796 16652
rect 11848 16640 11854 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 11848 16612 14105 16640
rect 11848 16600 11854 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 9858 16572 9864 16584
rect 4157 16535 4215 16541
rect 4264 16544 9864 16572
rect 3786 16464 3792 16516
rect 3844 16504 3850 16516
rect 4264 16504 4292 16544
rect 9858 16532 9864 16544
rect 9916 16532 9922 16584
rect 10042 16532 10048 16584
rect 10100 16532 10106 16584
rect 12802 16532 12808 16584
rect 12860 16532 12866 16584
rect 14274 16532 14280 16584
rect 14332 16532 14338 16584
rect 17310 16572 17316 16584
rect 16776 16544 17316 16572
rect 11054 16504 11060 16516
rect 3844 16476 4292 16504
rect 4632 16476 11060 16504
rect 3844 16464 3850 16476
rect 4632 16445 4660 16476
rect 11054 16464 11060 16476
rect 11112 16464 11118 16516
rect 12986 16464 12992 16516
rect 13044 16504 13050 16516
rect 16776 16513 16804 16544
rect 17310 16532 17316 16544
rect 17368 16532 17374 16584
rect 16761 16507 16819 16513
rect 16761 16504 16773 16507
rect 13044 16476 16773 16504
rect 13044 16464 13050 16476
rect 16761 16473 16773 16476
rect 16807 16473 16819 16507
rect 16761 16467 16819 16473
rect 16850 16464 16856 16516
rect 16908 16504 16914 16516
rect 18141 16507 18199 16513
rect 18141 16504 18153 16507
rect 16908 16476 18153 16504
rect 16908 16464 16914 16476
rect 18141 16473 18153 16476
rect 18187 16473 18199 16507
rect 18141 16467 18199 16473
rect 4617 16439 4675 16445
rect 4617 16405 4629 16439
rect 4663 16405 4675 16439
rect 4617 16399 4675 16405
rect 10137 16439 10195 16445
rect 10137 16405 10149 16439
rect 10183 16436 10195 16439
rect 10226 16436 10232 16448
rect 10183 16408 10232 16436
rect 10183 16405 10195 16408
rect 10137 16399 10195 16405
rect 10226 16396 10232 16408
rect 10284 16396 10290 16448
rect 12897 16439 12955 16445
rect 12897 16405 12909 16439
rect 12943 16436 12955 16439
rect 13630 16436 13636 16448
rect 12943 16408 13636 16436
rect 12943 16405 12955 16408
rect 12897 16399 12955 16405
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 16482 16396 16488 16448
rect 16540 16436 16546 16448
rect 16961 16439 17019 16445
rect 16961 16436 16973 16439
rect 16540 16408 16973 16436
rect 16540 16396 16546 16408
rect 16961 16405 16973 16408
rect 17007 16405 17019 16439
rect 16961 16399 17019 16405
rect 1104 16346 18860 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 7610 16346
rect 7662 16294 7674 16346
rect 7726 16294 7738 16346
rect 7790 16294 7802 16346
rect 7854 16294 7866 16346
rect 7918 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 17610 16346
rect 17662 16294 17674 16346
rect 17726 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 18860 16346
rect 1104 16272 18860 16294
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 3283 16204 9352 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 6914 16124 6920 16176
rect 6972 16164 6978 16176
rect 6972 16136 7696 16164
rect 6972 16124 6978 16136
rect 3050 16056 3056 16108
rect 3108 16096 3114 16108
rect 3145 16099 3203 16105
rect 3145 16096 3157 16099
rect 3108 16068 3157 16096
rect 3108 16056 3114 16068
rect 3145 16065 3157 16068
rect 3191 16065 3203 16099
rect 3145 16059 3203 16065
rect 3326 16056 3332 16108
rect 3384 16056 3390 16108
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 7668 16105 7696 16136
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 5684 16068 7481 16096
rect 5684 16056 5690 16068
rect 7469 16065 7481 16068
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 7653 16099 7711 16105
rect 7653 16065 7665 16099
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 9122 16056 9128 16108
rect 9180 16056 9186 16108
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 7340 16000 7757 16028
rect 7340 15988 7346 16000
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 8021 16031 8079 16037
rect 8021 16028 8033 16031
rect 7745 15991 7803 15997
rect 7852 16000 8033 16028
rect 2958 15920 2964 15972
rect 3016 15920 3022 15972
rect 4246 15920 4252 15972
rect 4304 15960 4310 15972
rect 7852 15960 7880 16000
rect 8021 15997 8033 16000
rect 8067 15997 8079 16031
rect 9324 16028 9352 16204
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 12802 16232 12808 16244
rect 9548 16204 12808 16232
rect 9548 16192 9554 16204
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 12894 16192 12900 16244
rect 12952 16192 12958 16244
rect 13004 16204 13492 16232
rect 9858 16124 9864 16176
rect 9916 16164 9922 16176
rect 13004 16164 13032 16204
rect 13464 16173 13492 16204
rect 14826 16192 14832 16244
rect 14884 16232 14890 16244
rect 14921 16235 14979 16241
rect 14921 16232 14933 16235
rect 14884 16204 14933 16232
rect 14884 16192 14890 16204
rect 14921 16201 14933 16204
rect 14967 16201 14979 16235
rect 14921 16195 14979 16201
rect 9916 16136 13032 16164
rect 13449 16167 13507 16173
rect 9916 16124 9922 16136
rect 13449 16133 13461 16167
rect 13495 16133 13507 16167
rect 16758 16164 16764 16176
rect 14674 16136 16764 16164
rect 13449 16127 13507 16133
rect 16758 16124 16764 16136
rect 16816 16124 16822 16176
rect 11146 16056 11152 16108
rect 11204 16096 11210 16108
rect 11204 16068 12756 16096
rect 11204 16056 11210 16068
rect 9324 16000 12572 16028
rect 8021 15991 8079 15997
rect 4304 15932 7880 15960
rect 12544 15960 12572 16000
rect 12618 15988 12624 16040
rect 12676 15988 12682 16040
rect 12728 16037 12756 16068
rect 15010 16056 15016 16108
rect 15068 16056 15074 16108
rect 15194 16056 15200 16108
rect 15252 16056 15258 16108
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 12713 16031 12771 16037
rect 12713 15997 12725 16031
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 12986 15988 12992 16040
rect 13044 15988 13050 16040
rect 13078 15988 13084 16040
rect 13136 15988 13142 16040
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 16028 13231 16031
rect 14090 16028 14096 16040
rect 13219 16000 14096 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 15488 16028 15516 16059
rect 14936 16000 15516 16028
rect 12802 15960 12808 15972
rect 12544 15932 12808 15960
rect 4304 15920 4310 15932
rect 12802 15920 12808 15932
rect 12860 15920 12866 15972
rect 3513 15895 3571 15901
rect 3513 15861 3525 15895
rect 3559 15892 3571 15895
rect 6822 15892 6828 15904
rect 3559 15864 6828 15892
rect 3559 15861 3571 15864
rect 3513 15855 3571 15861
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7466 15852 7472 15904
rect 7524 15852 7530 15904
rect 8018 15852 8024 15904
rect 8076 15892 8082 15904
rect 9493 15895 9551 15901
rect 9493 15892 9505 15895
rect 8076 15864 9505 15892
rect 8076 15852 8082 15864
rect 9493 15861 9505 15864
rect 9539 15861 9551 15895
rect 9493 15855 9551 15861
rect 12437 15895 12495 15901
rect 12437 15861 12449 15895
rect 12483 15892 12495 15895
rect 12526 15892 12532 15904
rect 12483 15864 12532 15892
rect 12483 15861 12495 15864
rect 12437 15855 12495 15861
rect 12526 15852 12532 15864
rect 12584 15852 12590 15904
rect 12820 15892 12848 15920
rect 13078 15892 13084 15904
rect 12820 15864 13084 15892
rect 13078 15852 13084 15864
rect 13136 15852 13142 15904
rect 13998 15852 14004 15904
rect 14056 15892 14062 15904
rect 14936 15892 14964 16000
rect 15764 15960 15792 16059
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16632 16068 16865 16096
rect 16632 16056 16638 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 18230 16056 18236 16108
rect 18288 16056 18294 16108
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 16028 17003 16031
rect 17494 16028 17500 16040
rect 16991 16000 17500 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17494 15988 17500 16000
rect 17552 15988 17558 16040
rect 18138 15960 18144 15972
rect 15764 15932 18144 15960
rect 18138 15920 18144 15932
rect 18196 15920 18202 15972
rect 14056 15864 14964 15892
rect 15013 15895 15071 15901
rect 14056 15852 14062 15864
rect 15013 15861 15025 15895
rect 15059 15892 15071 15895
rect 15102 15892 15108 15904
rect 15059 15864 15108 15892
rect 15059 15861 15071 15864
rect 15013 15855 15071 15861
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 15565 15895 15623 15901
rect 15565 15861 15577 15895
rect 15611 15892 15623 15895
rect 15746 15892 15752 15904
rect 15611 15864 15752 15892
rect 15611 15861 15623 15864
rect 15565 15855 15623 15861
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 15841 15895 15899 15901
rect 15841 15861 15853 15895
rect 15887 15892 15899 15895
rect 16574 15892 16580 15904
rect 15887 15864 16580 15892
rect 15887 15861 15899 15864
rect 15841 15855 15899 15861
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 17221 15895 17279 15901
rect 17221 15861 17233 15895
rect 17267 15892 17279 15895
rect 17402 15892 17408 15904
rect 17267 15864 17408 15892
rect 17267 15861 17279 15864
rect 17221 15855 17279 15861
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 18046 15852 18052 15904
rect 18104 15892 18110 15904
rect 18417 15895 18475 15901
rect 18417 15892 18429 15895
rect 18104 15864 18429 15892
rect 18104 15852 18110 15864
rect 18417 15861 18429 15864
rect 18463 15861 18475 15895
rect 18417 15855 18475 15861
rect 1104 15802 18860 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 16950 15802
rect 17002 15750 17014 15802
rect 17066 15750 17078 15802
rect 17130 15750 17142 15802
rect 17194 15750 17206 15802
rect 17258 15750 18860 15802
rect 1104 15728 18860 15750
rect 4985 15691 5043 15697
rect 4985 15657 4997 15691
rect 5031 15688 5043 15691
rect 8754 15688 8760 15700
rect 5031 15660 8760 15688
rect 5031 15657 5043 15660
rect 4985 15651 5043 15657
rect 8754 15648 8760 15660
rect 8812 15688 8818 15700
rect 9582 15688 9588 15700
rect 8812 15660 9588 15688
rect 8812 15648 8818 15660
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 11974 15688 11980 15700
rect 10796 15660 11980 15688
rect 10134 15620 10140 15632
rect 5000 15592 10140 15620
rect 5000 15564 5028 15592
rect 10134 15580 10140 15592
rect 10192 15620 10198 15632
rect 10796 15620 10824 15660
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 13170 15648 13176 15700
rect 13228 15688 13234 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 13228 15660 13461 15688
rect 13228 15648 13234 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 16850 15688 16856 15700
rect 13449 15651 13507 15657
rect 13556 15660 16856 15688
rect 12250 15620 12256 15632
rect 10192 15592 10824 15620
rect 11992 15592 12256 15620
rect 10192 15580 10198 15592
rect 4522 15512 4528 15564
rect 4580 15512 4586 15564
rect 4982 15512 4988 15564
rect 5040 15512 5046 15564
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 10594 15552 10600 15564
rect 6512 15524 10600 15552
rect 6512 15512 6518 15524
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 10689 15555 10747 15561
rect 10689 15521 10701 15555
rect 10735 15552 10747 15555
rect 11422 15552 11428 15564
rect 10735 15524 11428 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 11698 15512 11704 15564
rect 11756 15552 11762 15564
rect 11992 15552 12020 15592
rect 12250 15580 12256 15592
rect 12308 15580 12314 15632
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 13556 15620 13584 15660
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 12492 15592 13584 15620
rect 12492 15580 12498 15592
rect 11756 15524 12020 15552
rect 11756 15512 11762 15524
rect 12158 15512 12164 15564
rect 12216 15552 12222 15564
rect 15841 15555 15899 15561
rect 15841 15552 15853 15555
rect 12216 15524 15853 15552
rect 12216 15512 12222 15524
rect 15841 15521 15853 15524
rect 15887 15521 15899 15555
rect 15841 15515 15899 15521
rect 1489 15487 1547 15493
rect 1489 15453 1501 15487
rect 1535 15484 1547 15487
rect 5350 15484 5356 15496
rect 1535 15456 5356 15484
rect 1535 15453 1547 15456
rect 1489 15447 1547 15453
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 12308 15456 13645 15484
rect 12308 15444 12314 15456
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13906 15444 13912 15496
rect 13964 15444 13970 15496
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 3418 15376 3424 15428
rect 3476 15416 3482 15428
rect 3789 15419 3847 15425
rect 3789 15416 3801 15419
rect 3476 15388 3801 15416
rect 3476 15376 3482 15388
rect 3789 15385 3801 15388
rect 3835 15385 3847 15419
rect 3789 15379 3847 15385
rect 4801 15419 4859 15425
rect 4801 15385 4813 15419
rect 4847 15416 4859 15419
rect 10965 15419 11023 15425
rect 4847 15388 10778 15416
rect 4847 15385 4859 15388
rect 4801 15379 4859 15385
rect 1578 15308 1584 15360
rect 1636 15308 1642 15360
rect 4982 15308 4988 15360
rect 5040 15357 5046 15360
rect 5040 15351 5059 15357
rect 5047 15317 5059 15351
rect 5040 15311 5059 15317
rect 5040 15308 5046 15311
rect 5166 15308 5172 15360
rect 5224 15308 5230 15360
rect 8846 15308 8852 15360
rect 8904 15348 8910 15360
rect 9490 15348 9496 15360
rect 8904 15320 9496 15348
rect 8904 15308 8910 15320
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 10750 15348 10778 15388
rect 10965 15385 10977 15419
rect 11011 15416 11023 15419
rect 11238 15416 11244 15428
rect 11011 15388 11244 15416
rect 11011 15385 11023 15388
rect 10965 15379 11023 15385
rect 11238 15376 11244 15388
rect 11296 15376 11302 15428
rect 11348 15388 11454 15416
rect 12268 15388 13952 15416
rect 11348 15360 11376 15388
rect 11146 15348 11152 15360
rect 10750 15320 11152 15348
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 11330 15308 11336 15360
rect 11388 15308 11394 15360
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 12268 15348 12296 15388
rect 11756 15320 12296 15348
rect 11756 15308 11762 15320
rect 12802 15308 12808 15360
rect 12860 15348 12866 15360
rect 13722 15348 13728 15360
rect 12860 15320 13728 15348
rect 12860 15308 12866 15320
rect 13722 15308 13728 15320
rect 13780 15308 13786 15360
rect 13814 15308 13820 15360
rect 13872 15308 13878 15360
rect 13924 15348 13952 15388
rect 14366 15376 14372 15428
rect 14424 15376 14430 15428
rect 14476 15388 14858 15416
rect 14476 15348 14504 15388
rect 13924 15320 14504 15348
rect 1104 15258 18860 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 17610 15258
rect 17662 15206 17674 15258
rect 17726 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 18860 15258
rect 1104 15184 18860 15206
rect 10962 15104 10968 15156
rect 11020 15144 11026 15156
rect 11020 15116 11100 15144
rect 11020 15104 11026 15116
rect 6546 15036 6552 15088
rect 6604 15076 6610 15088
rect 10686 15076 10692 15088
rect 6604 15048 10692 15076
rect 6604 15036 6610 15048
rect 10686 15036 10692 15048
rect 10744 15036 10750 15088
rect 11072 15076 11100 15116
rect 11146 15104 11152 15156
rect 11204 15144 11210 15156
rect 11514 15144 11520 15156
rect 11204 15116 11520 15144
rect 11204 15104 11210 15116
rect 11514 15104 11520 15116
rect 11572 15144 11578 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 11572 15116 11805 15144
rect 11572 15104 11578 15116
rect 11793 15113 11805 15116
rect 11839 15113 11851 15147
rect 11793 15107 11851 15113
rect 11882 15104 11888 15156
rect 11940 15104 11946 15156
rect 11974 15104 11980 15156
rect 12032 15104 12038 15156
rect 12066 15104 12072 15156
rect 12124 15144 12130 15156
rect 12124 15116 17908 15144
rect 12124 15104 12130 15116
rect 11072 15048 11284 15076
rect 6086 14968 6092 15020
rect 6144 15008 6150 15020
rect 11146 15014 11152 15020
rect 11072 15008 11152 15014
rect 6144 14986 11152 15008
rect 6144 14980 11100 14986
rect 6144 14968 6150 14980
rect 11146 14968 11152 14986
rect 11204 14968 11210 15020
rect 11256 15017 11284 15048
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 15105 15079 15163 15085
rect 11664 15048 13110 15076
rect 11664 15036 11670 15048
rect 15105 15045 15117 15079
rect 15151 15076 15163 15079
rect 16298 15076 16304 15088
rect 15151 15048 16304 15076
rect 15151 15045 15163 15048
rect 15105 15039 15163 15045
rect 11241 15011 11299 15017
rect 11241 14977 11253 15011
rect 11287 14977 11299 15011
rect 11241 14971 11299 14977
rect 11422 14968 11428 15020
rect 11480 15008 11486 15020
rect 12342 15008 12348 15020
rect 11480 14980 12348 15008
rect 11480 14968 11486 14980
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 14734 14968 14740 15020
rect 14792 14968 14798 15020
rect 9582 14900 9588 14952
rect 9640 14940 9646 14952
rect 10778 14940 10784 14952
rect 9640 14912 10784 14940
rect 9640 14900 9646 14912
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 12621 14943 12679 14949
rect 11655 14912 12480 14940
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 6270 14832 6276 14884
rect 6328 14872 6334 14884
rect 12161 14875 12219 14881
rect 12161 14872 12173 14875
rect 6328 14844 12173 14872
rect 6328 14832 6334 14844
rect 12161 14841 12173 14844
rect 12207 14841 12219 14875
rect 12161 14835 12219 14841
rect 5074 14764 5080 14816
rect 5132 14804 5138 14816
rect 12066 14804 12072 14816
rect 5132 14776 12072 14804
rect 5132 14764 5138 14776
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 12452 14804 12480 14912
rect 12621 14909 12633 14943
rect 12667 14940 12679 14943
rect 12986 14940 12992 14952
rect 12667 14912 12992 14940
rect 12667 14909 12679 14912
rect 12621 14903 12679 14909
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 15120 14940 15148 15039
rect 16298 15036 16304 15048
rect 16356 15076 16362 15088
rect 16356 15048 17816 15076
rect 16356 15036 16362 15048
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15378 15008 15384 15020
rect 15243 14980 15384 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 17681 15011 17739 15017
rect 17681 15008 17693 15011
rect 17328 14980 17693 15008
rect 13136 14912 15148 14940
rect 13136 14900 13142 14912
rect 13906 14832 13912 14884
rect 13964 14872 13970 14884
rect 15102 14872 15108 14884
rect 13964 14844 15108 14872
rect 13964 14832 13970 14844
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 16942 14832 16948 14884
rect 17000 14872 17006 14884
rect 17328 14881 17356 14980
rect 17681 14977 17693 14980
rect 17727 14977 17739 15011
rect 17681 14971 17739 14977
rect 17788 14940 17816 15048
rect 17880 15017 17908 15116
rect 17865 15011 17923 15017
rect 17865 14977 17877 15011
rect 17911 14977 17923 15011
rect 17865 14971 17923 14977
rect 18690 14940 18696 14952
rect 17788 14912 18696 14940
rect 18690 14900 18696 14912
rect 18748 14900 18754 14952
rect 17313 14875 17371 14881
rect 17313 14872 17325 14875
rect 17000 14844 17325 14872
rect 17000 14832 17006 14844
rect 17313 14841 17325 14844
rect 17359 14841 17371 14875
rect 17313 14835 17371 14841
rect 13078 14804 13084 14816
rect 12452 14776 13084 14804
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 14093 14807 14151 14813
rect 14093 14804 14105 14807
rect 13412 14776 14105 14804
rect 13412 14764 13418 14776
rect 14093 14773 14105 14776
rect 14139 14773 14151 14807
rect 14093 14767 14151 14773
rect 15286 14764 15292 14816
rect 15344 14764 15350 14816
rect 16758 14764 16764 14816
rect 16816 14804 16822 14816
rect 17681 14807 17739 14813
rect 17681 14804 17693 14807
rect 16816 14776 17693 14804
rect 16816 14764 16822 14776
rect 17681 14773 17693 14776
rect 17727 14773 17739 14807
rect 17681 14767 17739 14773
rect 1104 14714 18860 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 16950 14714
rect 17002 14662 17014 14714
rect 17066 14662 17078 14714
rect 17130 14662 17142 14714
rect 17194 14662 17206 14714
rect 17258 14662 18860 14714
rect 1104 14640 18860 14662
rect 6546 14560 6552 14612
rect 6604 14560 6610 14612
rect 8386 14560 8392 14612
rect 8444 14600 8450 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 8444 14572 12265 14600
rect 8444 14560 8450 14572
rect 12253 14569 12265 14572
rect 12299 14600 12311 14603
rect 14734 14600 14740 14612
rect 12299 14572 14740 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 13906 14532 13912 14544
rect 3160 14504 13912 14532
rect 3160 14405 3188 14504
rect 13906 14492 13912 14504
rect 13964 14492 13970 14544
rect 14274 14492 14280 14544
rect 14332 14532 14338 14544
rect 17037 14535 17095 14541
rect 17037 14532 17049 14535
rect 14332 14504 17049 14532
rect 14332 14492 14338 14504
rect 17037 14501 17049 14504
rect 17083 14501 17095 14535
rect 17037 14495 17095 14501
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 11698 14464 11704 14476
rect 6319 14436 11704 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 11974 14464 11980 14476
rect 11931 14436 11980 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 15378 14464 15384 14476
rect 13596 14436 15384 14464
rect 13596 14424 13602 14436
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 16022 14424 16028 14476
rect 16080 14464 16086 14476
rect 17129 14467 17187 14473
rect 17129 14464 17141 14467
rect 16080 14436 17141 14464
rect 16080 14424 16086 14436
rect 17129 14433 17141 14436
rect 17175 14433 17187 14467
rect 17129 14427 17187 14433
rect 3145 14399 3203 14405
rect 3145 14365 3157 14399
rect 3191 14365 3203 14399
rect 3145 14359 3203 14365
rect 6086 14356 6092 14408
rect 6144 14396 6150 14408
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 6144 14368 6193 14396
rect 6144 14356 6150 14368
rect 6181 14365 6193 14368
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14396 6515 14399
rect 6546 14396 6552 14408
rect 6503 14368 6552 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 9398 14396 9404 14408
rect 6880 14368 9404 14396
rect 6880 14356 6886 14368
rect 9398 14356 9404 14368
rect 9456 14356 9462 14408
rect 11422 14356 11428 14408
rect 11480 14396 11486 14408
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11480 14368 11805 14396
rect 11480 14356 11486 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 13633 14399 13691 14405
rect 13633 14396 13645 14399
rect 11793 14359 11851 14365
rect 11900 14368 13645 14396
rect 2777 14331 2835 14337
rect 2777 14297 2789 14331
rect 2823 14328 2835 14331
rect 2866 14328 2872 14340
rect 2823 14300 2872 14328
rect 2823 14297 2835 14300
rect 2777 14291 2835 14297
rect 2866 14288 2872 14300
rect 2924 14328 2930 14340
rect 2924 14300 7052 14328
rect 2924 14288 2930 14300
rect 2958 14220 2964 14272
rect 3016 14220 3022 14272
rect 3050 14220 3056 14272
rect 3108 14220 3114 14272
rect 3329 14263 3387 14269
rect 3329 14229 3341 14263
rect 3375 14260 3387 14263
rect 6178 14260 6184 14272
rect 3375 14232 6184 14260
rect 3375 14229 3387 14232
rect 3329 14223 3387 14229
rect 6178 14220 6184 14232
rect 6236 14220 6242 14272
rect 7024 14260 7052 14300
rect 11606 14288 11612 14340
rect 11664 14328 11670 14340
rect 11900 14328 11928 14368
rect 13633 14365 13645 14368
rect 13679 14365 13691 14399
rect 13633 14359 13691 14365
rect 14826 14356 14832 14408
rect 14884 14396 14890 14408
rect 17037 14399 17095 14405
rect 17037 14396 17049 14399
rect 14884 14368 17049 14396
rect 14884 14356 14890 14368
rect 17037 14365 17049 14368
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 11664 14300 11928 14328
rect 12069 14331 12127 14337
rect 11664 14288 11670 14300
rect 12069 14297 12081 14331
rect 12115 14328 12127 14331
rect 14458 14328 14464 14340
rect 12115 14300 14464 14328
rect 12115 14297 12127 14300
rect 12069 14291 12127 14297
rect 12084 14260 12112 14291
rect 14458 14288 14464 14300
rect 14516 14288 14522 14340
rect 15194 14288 15200 14340
rect 15252 14328 15258 14340
rect 15654 14328 15660 14340
rect 15252 14300 15660 14328
rect 15252 14288 15258 14300
rect 15654 14288 15660 14300
rect 15712 14328 15718 14340
rect 17313 14331 17371 14337
rect 17313 14328 17325 14331
rect 15712 14300 17325 14328
rect 15712 14288 15718 14300
rect 17313 14297 17325 14300
rect 17359 14297 17371 14331
rect 17313 14291 17371 14297
rect 7024 14232 12112 14260
rect 12250 14220 12256 14272
rect 12308 14269 12314 14272
rect 12308 14263 12327 14269
rect 12315 14229 12327 14263
rect 12308 14223 12327 14229
rect 12308 14220 12314 14223
rect 12434 14220 12440 14272
rect 12492 14220 12498 14272
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14260 13507 14263
rect 15838 14260 15844 14272
rect 13495 14232 15844 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 1104 14170 18860 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 17610 14170
rect 17662 14118 17674 14170
rect 17726 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 18860 14170
rect 1104 14096 18860 14118
rect 3050 14016 3056 14068
rect 3108 14056 3114 14068
rect 14826 14056 14832 14068
rect 3108 14028 14832 14056
rect 3108 14016 3114 14028
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 4062 13988 4068 14000
rect 4002 13960 4068 13988
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 5902 13948 5908 14000
rect 5960 13988 5966 14000
rect 6546 13988 6552 14000
rect 5960 13960 6552 13988
rect 5960 13948 5966 13960
rect 6546 13948 6552 13960
rect 6604 13948 6610 14000
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 13538 13988 13544 14000
rect 11204 13960 13544 13988
rect 11204 13948 11210 13960
rect 13538 13948 13544 13960
rect 13596 13948 13602 14000
rect 2498 13880 2504 13932
rect 2556 13880 2562 13932
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13920 4491 13923
rect 5920 13920 5948 13948
rect 4479 13892 5948 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 6178 13880 6184 13932
rect 6236 13920 6242 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6236 13892 6837 13920
rect 6236 13880 6242 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 8570 13880 8576 13932
rect 8628 13880 8634 13932
rect 10870 13880 10876 13932
rect 10928 13920 10934 13932
rect 13170 13920 13176 13932
rect 10928 13892 13176 13920
rect 10928 13880 10934 13892
rect 13170 13880 13176 13892
rect 13228 13880 13234 13932
rect 15194 13880 15200 13932
rect 15252 13880 15258 13932
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13852 2283 13855
rect 2777 13855 2835 13861
rect 2777 13852 2789 13855
rect 2271 13824 2789 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 2777 13821 2789 13824
rect 2823 13852 2835 13855
rect 3510 13852 3516 13864
rect 2823 13824 3516 13852
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 4338 13852 4344 13864
rect 4295 13824 4344 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 4338 13812 4344 13824
rect 4396 13812 4402 13864
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 5718 13852 5724 13864
rect 4571 13824 5724 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 6546 13852 6552 13864
rect 6420 13824 6552 13852
rect 6420 13812 6426 13824
rect 6546 13812 6552 13824
rect 6604 13852 6610 13864
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 6604 13824 7205 13852
rect 6604 13812 6610 13824
rect 7193 13821 7205 13824
rect 7239 13821 7251 13855
rect 7469 13855 7527 13861
rect 7469 13852 7481 13855
rect 7193 13815 7251 13821
rect 7300 13824 7481 13852
rect 4154 13744 4160 13796
rect 4212 13784 4218 13796
rect 7300 13784 7328 13824
rect 7469 13821 7481 13824
rect 7515 13821 7527 13855
rect 7469 13815 7527 13821
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8941 13855 8999 13861
rect 8941 13852 8953 13855
rect 8536 13824 8953 13852
rect 8536 13812 8542 13824
rect 8941 13821 8953 13824
rect 8987 13821 8999 13855
rect 8941 13815 8999 13821
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 11422 13852 11428 13864
rect 11204 13824 11428 13852
rect 11204 13812 11210 13824
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 12216 13824 13829 13852
rect 12216 13812 12222 13824
rect 13817 13821 13829 13824
rect 13863 13852 13875 13855
rect 14182 13852 14188 13864
rect 13863 13824 14188 13852
rect 13863 13821 13875 13824
rect 13817 13815 13875 13821
rect 14182 13812 14188 13824
rect 14240 13812 14246 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13852 15623 13855
rect 16114 13852 16120 13864
rect 15611 13824 16120 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 16114 13812 16120 13824
rect 16172 13812 16178 13864
rect 4212 13756 7328 13784
rect 4212 13744 4218 13756
rect 4890 13676 4896 13728
rect 4948 13716 4954 13728
rect 6914 13716 6920 13728
rect 4948 13688 6920 13716
rect 4948 13676 4954 13688
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 7009 13719 7067 13725
rect 7009 13685 7021 13719
rect 7055 13716 7067 13719
rect 7282 13716 7288 13728
rect 7055 13688 7288 13716
rect 7055 13685 7067 13688
rect 7009 13679 7067 13685
rect 7282 13676 7288 13688
rect 7340 13716 7346 13728
rect 9030 13716 9036 13728
rect 7340 13688 9036 13716
rect 7340 13676 7346 13688
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13538 13716 13544 13728
rect 13136 13688 13544 13716
rect 13136 13676 13142 13688
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 14080 13719 14138 13725
rect 14080 13685 14092 13719
rect 14126 13716 14138 13719
rect 15470 13716 15476 13728
rect 14126 13688 15476 13716
rect 14126 13685 14138 13688
rect 14080 13679 14138 13685
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 1104 13626 18860 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 16950 13626
rect 17002 13574 17014 13626
rect 17066 13574 17078 13626
rect 17130 13574 17142 13626
rect 17194 13574 17206 13626
rect 17258 13574 18860 13626
rect 1104 13552 18860 13574
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 6914 13512 6920 13524
rect 4580 13484 6920 13512
rect 4580 13472 4586 13484
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7466 13472 7472 13524
rect 7524 13472 7530 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 17313 13515 17371 13521
rect 17313 13512 17325 13515
rect 13320 13484 17325 13512
rect 13320 13472 13326 13484
rect 17313 13481 17325 13484
rect 17359 13481 17371 13515
rect 17313 13475 17371 13481
rect 4430 13404 4436 13456
rect 4488 13444 4494 13456
rect 7484 13444 7512 13472
rect 10594 13444 10600 13456
rect 4488 13416 10600 13444
rect 4488 13404 4494 13416
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 10962 13404 10968 13456
rect 11020 13444 11026 13456
rect 13078 13444 13084 13456
rect 11020 13416 13084 13444
rect 11020 13404 11026 13416
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 14918 13404 14924 13456
rect 14976 13444 14982 13456
rect 15289 13447 15347 13453
rect 15289 13444 15301 13447
rect 14976 13416 15301 13444
rect 14976 13404 14982 13416
rect 15289 13413 15301 13416
rect 15335 13413 15347 13447
rect 15289 13407 15347 13413
rect 7466 13376 7472 13388
rect 2976 13348 7472 13376
rect 2130 13268 2136 13320
rect 2188 13268 2194 13320
rect 2406 13268 2412 13320
rect 2464 13268 2470 13320
rect 2976 13317 3004 13348
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 8110 13336 8116 13388
rect 8168 13376 8174 13388
rect 8168 13348 15148 13376
rect 8168 13336 8174 13348
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13277 2651 13311
rect 2593 13271 2651 13277
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13277 3019 13311
rect 2961 13271 3019 13277
rect 2314 13200 2320 13252
rect 2372 13200 2378 13252
rect 2608 13240 2636 13271
rect 3142 13268 3148 13320
rect 3200 13268 3206 13320
rect 3789 13311 3847 13317
rect 3789 13277 3801 13311
rect 3835 13308 3847 13311
rect 4522 13308 4528 13320
rect 3835 13280 4528 13308
rect 3835 13277 3847 13280
rect 3789 13271 3847 13277
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 5534 13268 5540 13320
rect 5592 13308 5598 13320
rect 6086 13308 6092 13320
rect 5592 13280 6092 13308
rect 5592 13268 5598 13280
rect 6086 13268 6092 13280
rect 6144 13308 6150 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6144 13280 6285 13308
rect 6144 13268 6150 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 7098 13268 7104 13320
rect 7156 13308 7162 13320
rect 8938 13308 8944 13320
rect 7156 13280 8944 13308
rect 7156 13268 7162 13280
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 10042 13268 10048 13320
rect 10100 13308 10106 13320
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 10100 13280 10609 13308
rect 10100 13268 10106 13280
rect 10597 13277 10609 13280
rect 10643 13308 10655 13311
rect 10870 13308 10876 13320
rect 10643 13280 10876 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13504 13280 13737 13308
rect 13504 13268 13510 13280
rect 13725 13277 13737 13280
rect 13771 13308 13783 13311
rect 13998 13308 14004 13320
rect 13771 13280 14004 13308
rect 13771 13277 13783 13280
rect 13725 13271 13783 13277
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13308 14519 13311
rect 14734 13308 14740 13320
rect 14507 13280 14740 13308
rect 14507 13277 14519 13280
rect 14461 13271 14519 13277
rect 14734 13268 14740 13280
rect 14792 13268 14798 13320
rect 15120 13317 15148 13348
rect 15838 13336 15844 13388
rect 15896 13336 15902 13388
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13277 15163 13311
rect 15105 13271 15163 13277
rect 15562 13268 15568 13320
rect 15620 13268 15626 13320
rect 3510 13240 3516 13252
rect 2608 13212 3516 13240
rect 3510 13200 3516 13212
rect 3568 13200 3574 13252
rect 13814 13200 13820 13252
rect 13872 13200 13878 13252
rect 14090 13200 14096 13252
rect 14148 13200 14154 13252
rect 16298 13200 16304 13252
rect 16356 13200 16362 13252
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 5994 13172 6000 13184
rect 3927 13144 6000 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 5994 13132 6000 13144
rect 6052 13132 6058 13184
rect 6362 13132 6368 13184
rect 6420 13132 6426 13184
rect 6638 13132 6644 13184
rect 6696 13172 6702 13184
rect 9582 13172 9588 13184
rect 6696 13144 9588 13172
rect 6696 13132 6702 13144
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 10686 13132 10692 13184
rect 10744 13132 10750 13184
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 14277 13175 14335 13181
rect 14277 13172 14289 13175
rect 11940 13144 14289 13172
rect 11940 13132 11946 13144
rect 14277 13141 14289 13144
rect 14323 13141 14335 13175
rect 14277 13135 14335 13141
rect 14369 13175 14427 13181
rect 14369 13141 14381 13175
rect 14415 13172 14427 13175
rect 14458 13172 14464 13184
rect 14415 13144 14464 13172
rect 14415 13141 14427 13144
rect 14369 13135 14427 13141
rect 14458 13132 14464 13144
rect 14516 13132 14522 13184
rect 14642 13132 14648 13184
rect 14700 13132 14706 13184
rect 1104 13082 18860 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 17610 13082
rect 17662 13030 17674 13082
rect 17726 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 18860 13082
rect 1104 13008 18860 13030
rect 1397 12971 1455 12977
rect 1397 12937 1409 12971
rect 1443 12968 1455 12971
rect 5626 12968 5632 12980
rect 1443 12940 5632 12968
rect 1443 12937 1455 12940
rect 1397 12931 1455 12937
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 10134 12968 10140 12980
rect 7616 12940 10140 12968
rect 7616 12928 7622 12940
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11606 12968 11612 12980
rect 11020 12940 11612 12968
rect 11020 12928 11026 12940
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12250 12928 12256 12980
rect 12308 12968 12314 12980
rect 13262 12968 13268 12980
rect 12308 12940 13268 12968
rect 12308 12928 12314 12940
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 14918 12928 14924 12980
rect 14976 12968 14982 12980
rect 16298 12968 16304 12980
rect 14976 12940 16304 12968
rect 14976 12928 14982 12940
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18233 12971 18291 12977
rect 18233 12968 18245 12971
rect 18196 12940 18245 12968
rect 18196 12928 18202 12940
rect 18233 12937 18245 12940
rect 18279 12968 18291 12971
rect 18414 12968 18420 12980
rect 18279 12940 18420 12968
rect 18279 12937 18291 12940
rect 18233 12931 18291 12937
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 5534 12900 5540 12912
rect 4094 12872 5540 12900
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 6546 12860 6552 12912
rect 6604 12900 6610 12912
rect 6604 12872 7696 12900
rect 6604 12860 6610 12872
rect 1578 12792 1584 12844
rect 1636 12792 1642 12844
rect 6178 12792 6184 12844
rect 6236 12832 6242 12844
rect 6638 12832 6644 12844
rect 6236 12804 6644 12832
rect 6236 12792 6242 12804
rect 6638 12792 6644 12804
rect 6696 12832 6702 12844
rect 7668 12841 7696 12872
rect 7834 12860 7840 12912
rect 7892 12900 7898 12912
rect 7892 12872 8418 12900
rect 7892 12860 7898 12872
rect 10686 12860 10692 12912
rect 10744 12900 10750 12912
rect 10744 12872 15502 12900
rect 10744 12860 10750 12872
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 6696 12804 7205 12832
rect 6696 12792 6702 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 2593 12767 2651 12773
rect 2593 12733 2605 12767
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12764 2927 12767
rect 7098 12764 7104 12776
rect 2915 12736 7104 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 2608 12628 2636 12727
rect 7098 12724 7104 12736
rect 7156 12724 7162 12776
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12764 7343 12767
rect 7558 12764 7564 12776
rect 7331 12736 7564 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 7558 12724 7564 12736
rect 7616 12724 7622 12776
rect 7668 12764 7696 12795
rect 18138 12792 18144 12844
rect 18196 12792 18202 12844
rect 7929 12767 7987 12773
rect 7668 12736 7788 12764
rect 3878 12656 3884 12708
rect 3936 12696 3942 12708
rect 4154 12696 4160 12708
rect 3936 12668 4160 12696
rect 3936 12656 3942 12668
rect 4154 12656 4160 12668
rect 4212 12656 4218 12708
rect 4890 12696 4896 12708
rect 4264 12668 4896 12696
rect 4264 12628 4292 12668
rect 4890 12656 4896 12668
rect 4948 12656 4954 12708
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 7650 12696 7656 12708
rect 5684 12668 7656 12696
rect 5684 12656 5690 12668
rect 7650 12656 7656 12668
rect 7708 12656 7714 12708
rect 7760 12640 7788 12736
rect 7929 12733 7941 12767
rect 7975 12764 7987 12767
rect 9122 12764 9128 12776
rect 7975 12736 9128 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 9122 12724 9128 12736
rect 9180 12724 9186 12776
rect 9214 12724 9220 12776
rect 9272 12764 9278 12776
rect 9401 12767 9459 12773
rect 9401 12764 9413 12767
rect 9272 12736 9413 12764
rect 9272 12724 9278 12736
rect 9401 12733 9413 12736
rect 9447 12764 9459 12767
rect 11422 12764 11428 12776
rect 9447 12736 11428 12764
rect 9447 12733 9459 12736
rect 9401 12727 9459 12733
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 11514 12724 11520 12776
rect 11572 12764 11578 12776
rect 11698 12764 11704 12776
rect 11572 12736 11704 12764
rect 11572 12724 11578 12736
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 14734 12764 14740 12776
rect 14240 12736 14740 12764
rect 14240 12724 14246 12736
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14844 12736 15025 12764
rect 9490 12656 9496 12708
rect 9548 12696 9554 12708
rect 14844 12696 14872 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 16574 12764 16580 12776
rect 16264 12736 16580 12764
rect 16264 12724 16270 12736
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 9548 12668 14872 12696
rect 9548 12656 9554 12668
rect 16390 12656 16396 12708
rect 16448 12696 16454 12708
rect 16448 12668 16896 12696
rect 16448 12656 16454 12668
rect 16868 12640 16896 12668
rect 2608 12600 4292 12628
rect 4338 12588 4344 12640
rect 4396 12588 4402 12640
rect 4706 12588 4712 12640
rect 4764 12628 4770 12640
rect 7561 12631 7619 12637
rect 7561 12628 7573 12631
rect 4764 12600 7573 12628
rect 4764 12588 4770 12600
rect 7561 12597 7573 12600
rect 7607 12597 7619 12631
rect 7561 12591 7619 12597
rect 7742 12588 7748 12640
rect 7800 12588 7806 12640
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 15102 12628 15108 12640
rect 14424 12600 15108 12628
rect 14424 12588 14430 12600
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 16485 12631 16543 12637
rect 16485 12597 16497 12631
rect 16531 12628 16543 12631
rect 16758 12628 16764 12640
rect 16531 12600 16764 12628
rect 16531 12597 16543 12600
rect 16485 12591 16543 12597
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 16850 12588 16856 12640
rect 16908 12588 16914 12640
rect 1104 12538 18860 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 16950 12538
rect 17002 12486 17014 12538
rect 17066 12486 17078 12538
rect 17130 12486 17142 12538
rect 17194 12486 17206 12538
rect 17258 12486 18860 12538
rect 1104 12464 18860 12486
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 3878 12424 3884 12436
rect 2087 12396 3884 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 4396 12396 8892 12424
rect 4396 12384 4402 12396
rect 2961 12359 3019 12365
rect 2961 12325 2973 12359
rect 3007 12356 3019 12359
rect 4246 12356 4252 12368
rect 3007 12328 4252 12356
rect 3007 12325 3019 12328
rect 2961 12319 3019 12325
rect 4246 12316 4252 12328
rect 4304 12316 4310 12368
rect 4890 12316 4896 12368
rect 4948 12356 4954 12368
rect 8386 12356 8392 12368
rect 4948 12328 8392 12356
rect 4948 12316 4954 12328
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 8864 12356 8892 12396
rect 8938 12384 8944 12436
rect 8996 12384 9002 12436
rect 9953 12427 10011 12433
rect 9953 12393 9965 12427
rect 9999 12424 10011 12427
rect 10042 12424 10048 12436
rect 9999 12396 10048 12424
rect 9999 12393 10011 12396
rect 9953 12387 10011 12393
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 10594 12384 10600 12436
rect 10652 12424 10658 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10652 12396 10701 12424
rect 10652 12384 10658 12396
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 10689 12387 10747 12393
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 11756 12396 14473 12424
rect 11756 12384 11762 12396
rect 14461 12393 14473 12396
rect 14507 12393 14519 12427
rect 14461 12387 14519 12393
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 16758 12424 16764 12436
rect 16632 12396 16764 12424
rect 16632 12384 16638 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 8864 12328 9444 12356
rect 3050 12288 3056 12300
rect 2240 12260 3056 12288
rect 2240 12229 2268 12260
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 3237 12291 3295 12297
rect 3237 12257 3249 12291
rect 3283 12288 3295 12291
rect 5258 12288 5264 12300
rect 3283 12260 5264 12288
rect 3283 12257 3295 12260
rect 3237 12251 3295 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 6270 12248 6276 12300
rect 6328 12248 6334 12300
rect 6362 12248 6368 12300
rect 6420 12248 6426 12300
rect 6546 12248 6552 12300
rect 6604 12248 6610 12300
rect 8294 12248 8300 12300
rect 8352 12288 8358 12300
rect 9416 12297 9444 12328
rect 10870 12316 10876 12368
rect 10928 12316 10934 12368
rect 14274 12356 14280 12368
rect 11624 12328 14280 12356
rect 9217 12291 9275 12297
rect 9217 12288 9229 12291
rect 8352 12260 9229 12288
rect 8352 12248 8358 12260
rect 9217 12257 9229 12260
rect 9263 12257 9275 12291
rect 9217 12251 9275 12257
rect 9401 12291 9459 12297
rect 9401 12257 9413 12291
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 9582 12248 9588 12300
rect 9640 12248 9646 12300
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12220 2559 12223
rect 2866 12220 2872 12232
rect 2547 12192 2872 12220
rect 2547 12189 2559 12192
rect 2501 12183 2559 12189
rect 2866 12180 2872 12192
rect 2924 12220 2930 12232
rect 3436 12229 3556 12230
rect 3145 12223 3203 12229
rect 3145 12220 3157 12223
rect 2924 12192 3157 12220
rect 2924 12180 2930 12192
rect 3145 12189 3157 12192
rect 3191 12189 3203 12223
rect 3145 12183 3203 12189
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3421 12223 3556 12229
rect 3421 12189 3433 12223
rect 3467 12202 3556 12223
rect 3467 12189 3479 12202
rect 3421 12183 3479 12189
rect 2409 12087 2467 12093
rect 2409 12053 2421 12087
rect 2455 12084 2467 12087
rect 2498 12084 2504 12096
rect 2455 12056 2504 12084
rect 2455 12053 2467 12056
rect 2409 12047 2467 12053
rect 2498 12044 2504 12056
rect 2556 12044 2562 12096
rect 3344 12084 3372 12183
rect 3528 12152 3556 12202
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 4120 12192 6469 12220
rect 4120 12180 4126 12192
rect 6457 12189 6469 12192
rect 6503 12220 6515 12223
rect 6638 12220 6644 12232
rect 6503 12192 6644 12220
rect 6503 12189 6515 12192
rect 6457 12183 6515 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6972 12192 7297 12220
rect 6972 12180 6978 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 9088 12192 9137 12220
rect 9088 12180 9094 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9674 12220 9680 12232
rect 9355 12192 9680 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12220 9827 12223
rect 9858 12220 9864 12232
rect 9815 12192 9864 12220
rect 9815 12189 9827 12192
rect 9769 12183 9827 12189
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 11624 12220 11652 12328
rect 14274 12316 14280 12328
rect 14332 12316 14338 12368
rect 16298 12316 16304 12368
rect 16356 12356 16362 12368
rect 17310 12356 17316 12368
rect 16356 12328 17316 12356
rect 16356 12316 16362 12328
rect 17310 12316 17316 12328
rect 17368 12316 17374 12368
rect 13722 12248 13728 12300
rect 13780 12288 13786 12300
rect 14550 12288 14556 12300
rect 13780 12260 14556 12288
rect 13780 12248 13786 12260
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 10336 12192 11652 12220
rect 7098 12152 7104 12164
rect 3528 12124 7104 12152
rect 7098 12112 7104 12124
rect 7156 12152 7162 12164
rect 8018 12152 8024 12164
rect 7156 12124 8024 12152
rect 7156 12112 7162 12124
rect 8018 12112 8024 12124
rect 8076 12112 8082 12164
rect 8478 12112 8484 12164
rect 8536 12152 8542 12164
rect 10336 12161 10364 12192
rect 14090 12180 14096 12232
rect 14148 12180 14154 12232
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 10321 12155 10379 12161
rect 10321 12152 10333 12155
rect 8536 12124 10333 12152
rect 8536 12112 8542 12124
rect 10321 12121 10333 12124
rect 10367 12121 10379 12155
rect 10321 12115 10379 12121
rect 10410 12112 10416 12164
rect 10468 12152 10474 12164
rect 11790 12152 11796 12164
rect 10468 12124 11796 12152
rect 10468 12112 10474 12124
rect 11790 12112 11796 12124
rect 11848 12112 11854 12164
rect 13446 12112 13452 12164
rect 13504 12152 13510 12164
rect 13722 12152 13728 12164
rect 13504 12124 13728 12152
rect 13504 12112 13510 12124
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 5074 12084 5080 12096
rect 3344 12056 5080 12084
rect 5074 12044 5080 12056
rect 5132 12044 5138 12096
rect 6086 12044 6092 12096
rect 6144 12044 6150 12096
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 6972 12056 7389 12084
rect 6972 12044 6978 12056
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 7377 12047 7435 12053
rect 9582 12044 9588 12096
rect 9640 12084 9646 12096
rect 10226 12084 10232 12096
rect 9640 12056 10232 12084
rect 9640 12044 9646 12056
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10686 12044 10692 12096
rect 10744 12093 10750 12096
rect 10744 12047 10756 12093
rect 10744 12044 10750 12047
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 11514 12084 11520 12096
rect 11388 12056 11520 12084
rect 11388 12044 11394 12056
rect 11514 12044 11520 12056
rect 11572 12044 11578 12096
rect 11882 12044 11888 12096
rect 11940 12084 11946 12096
rect 15838 12084 15844 12096
rect 11940 12056 15844 12084
rect 11940 12044 11946 12056
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 1104 11994 18860 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 17610 11994
rect 17662 11942 17674 11994
rect 17726 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 18860 11994
rect 1104 11920 18860 11942
rect 3326 11840 3332 11892
rect 3384 11880 3390 11892
rect 3878 11880 3884 11892
rect 3384 11852 3884 11880
rect 3384 11840 3390 11852
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 6365 11883 6423 11889
rect 6365 11849 6377 11883
rect 6411 11880 6423 11883
rect 6730 11880 6736 11892
rect 6411 11852 6736 11880
rect 6411 11849 6423 11852
rect 6365 11843 6423 11849
rect 6730 11840 6736 11852
rect 6788 11840 6794 11892
rect 9674 11880 9680 11892
rect 6932 11852 9680 11880
rect 5166 11812 5172 11824
rect 2148 11784 5172 11812
rect 1946 11704 1952 11756
rect 2004 11704 2010 11756
rect 2148 11753 2176 11784
rect 5166 11772 5172 11784
rect 5224 11772 5230 11824
rect 5276 11784 6684 11812
rect 2133 11747 2191 11753
rect 2133 11713 2145 11747
rect 2179 11713 2191 11747
rect 2133 11707 2191 11713
rect 2314 11704 2320 11756
rect 2372 11704 2378 11756
rect 2498 11704 2504 11756
rect 2556 11744 2562 11756
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2556 11716 2605 11744
rect 2556 11704 2562 11716
rect 2593 11713 2605 11716
rect 2639 11713 2651 11747
rect 2786 11747 2844 11753
rect 2786 11744 2798 11747
rect 2593 11707 2651 11713
rect 2700 11716 2798 11744
rect 1854 11568 1860 11620
rect 1912 11608 1918 11620
rect 2700 11608 2728 11716
rect 2786 11713 2798 11716
rect 2832 11713 2844 11747
rect 2786 11707 2844 11713
rect 3050 11704 3056 11756
rect 3108 11744 3114 11756
rect 3326 11744 3332 11756
rect 3108 11716 3332 11744
rect 3108 11704 3114 11716
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 4614 11704 4620 11756
rect 4672 11744 4678 11756
rect 5276 11744 5304 11784
rect 6656 11753 6684 11784
rect 4672 11716 5304 11744
rect 6641 11747 6699 11753
rect 4672 11704 4678 11716
rect 6641 11713 6653 11747
rect 6687 11713 6699 11747
rect 6932 11744 6960 11852
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 10410 11840 10416 11892
rect 10468 11840 10474 11892
rect 11790 11840 11796 11892
rect 11848 11880 11854 11892
rect 13446 11880 13452 11892
rect 11848 11852 13452 11880
rect 11848 11840 11854 11852
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 14001 11883 14059 11889
rect 14001 11849 14013 11883
rect 14047 11880 14059 11883
rect 14090 11880 14096 11892
rect 14047 11852 14096 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 9030 11772 9036 11824
rect 9088 11812 9094 11824
rect 10428 11812 10456 11840
rect 9088 11784 10456 11812
rect 9088 11772 9094 11784
rect 13170 11772 13176 11824
rect 13228 11772 13234 11824
rect 6641 11707 6699 11713
rect 6748 11716 6960 11744
rect 7009 11747 7067 11753
rect 6748 11688 6776 11716
rect 7009 11713 7021 11747
rect 7055 11744 7067 11747
rect 8110 11744 8116 11756
rect 7055 11716 8116 11744
rect 7055 11713 7067 11716
rect 7009 11707 7067 11713
rect 8110 11704 8116 11716
rect 8168 11704 8174 11756
rect 10410 11753 10416 11756
rect 10409 11707 10416 11753
rect 10468 11744 10474 11756
rect 11882 11744 11888 11756
rect 10468 11716 10509 11744
rect 11716 11716 11888 11744
rect 10410 11704 10416 11707
rect 10468 11704 10474 11716
rect 2958 11636 2964 11688
rect 3016 11676 3022 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 3016 11648 3433 11676
rect 3016 11636 3022 11648
rect 3421 11645 3433 11648
rect 3467 11676 3479 11679
rect 4890 11676 4896 11688
rect 3467 11648 4896 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 6362 11636 6368 11688
rect 6420 11636 6426 11688
rect 6546 11636 6552 11688
rect 6604 11636 6610 11688
rect 6730 11636 6736 11688
rect 6788 11636 6794 11688
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 8662 11676 8668 11688
rect 6871 11648 8668 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 1912 11580 2728 11608
rect 1912 11568 1918 11580
rect 4246 11568 4252 11620
rect 4304 11608 4310 11620
rect 6380 11608 6408 11636
rect 4304 11580 6408 11608
rect 4304 11568 4310 11580
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 7024 11540 7052 11648
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 10505 11679 10563 11685
rect 10505 11676 10517 11679
rect 9968 11648 10517 11676
rect 9968 11620 9996 11648
rect 10505 11645 10517 11648
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 10594 11636 10600 11688
rect 10652 11636 10658 11688
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11676 10747 11679
rect 11716 11676 11744 11716
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 15562 11744 15568 11756
rect 14231 11716 15568 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 10735 11648 11744 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 11848 11648 12265 11676
rect 11848 11636 11854 11648
rect 12253 11645 12265 11648
rect 12299 11676 12311 11679
rect 14200 11676 14228 11707
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 12299 11648 14228 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 7466 11568 7472 11620
rect 7524 11568 7530 11620
rect 7650 11568 7656 11620
rect 7708 11608 7714 11620
rect 9950 11608 9956 11620
rect 7708 11580 9956 11608
rect 7708 11568 7714 11580
rect 9950 11568 9956 11580
rect 10008 11568 10014 11620
rect 10152 11580 10456 11608
rect 6420 11512 7052 11540
rect 6420 11500 6426 11512
rect 7098 11500 7104 11552
rect 7156 11500 7162 11552
rect 8662 11500 8668 11552
rect 8720 11540 8726 11552
rect 10152 11540 10180 11580
rect 8720 11512 10180 11540
rect 10229 11543 10287 11549
rect 8720 11500 8726 11512
rect 10229 11509 10241 11543
rect 10275 11540 10287 11543
rect 10318 11540 10324 11552
rect 10275 11512 10324 11540
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 10428 11540 10456 11580
rect 11698 11540 11704 11552
rect 10428 11512 11704 11540
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12516 11543 12574 11549
rect 12516 11509 12528 11543
rect 12562 11540 12574 11543
rect 12986 11540 12992 11552
rect 12562 11512 12992 11540
rect 12562 11509 12574 11512
rect 12516 11503 12574 11509
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 14369 11543 14427 11549
rect 14369 11540 14381 11543
rect 14148 11512 14381 11540
rect 14148 11500 14154 11512
rect 14369 11509 14381 11512
rect 14415 11540 14427 11543
rect 14734 11540 14740 11552
rect 14415 11512 14740 11540
rect 14415 11509 14427 11512
rect 14369 11503 14427 11509
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 18138 11540 18144 11552
rect 17276 11512 18144 11540
rect 17276 11500 17282 11512
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 1104 11450 18860 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 16950 11450
rect 17002 11398 17014 11450
rect 17066 11398 17078 11450
rect 17130 11398 17142 11450
rect 17194 11398 17206 11450
rect 17258 11398 18860 11450
rect 1104 11376 18860 11398
rect 3786 11296 3792 11348
rect 3844 11296 3850 11348
rect 4522 11296 4528 11348
rect 4580 11296 4586 11348
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 8662 11336 8668 11348
rect 5868 11308 8668 11336
rect 5868 11296 5874 11308
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 8941 11339 8999 11345
rect 8941 11305 8953 11339
rect 8987 11336 8999 11339
rect 9122 11336 9128 11348
rect 8987 11308 9128 11336
rect 8987 11305 8999 11308
rect 8941 11299 8999 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10778 11336 10784 11348
rect 10652 11308 10784 11336
rect 10652 11296 10658 11308
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11112 11308 12388 11336
rect 11112 11296 11118 11308
rect 6546 11268 6552 11280
rect 4816 11240 6552 11268
rect 4062 11160 4068 11212
rect 4120 11160 4126 11212
rect 4430 11160 4436 11212
rect 4488 11160 4494 11212
rect 4816 11209 4844 11240
rect 6546 11228 6552 11240
rect 6604 11228 6610 11280
rect 9398 11228 9404 11280
rect 9456 11268 9462 11280
rect 9953 11271 10011 11277
rect 9456 11240 9904 11268
rect 9456 11228 9462 11240
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11169 4859 11203
rect 4801 11163 4859 11169
rect 4893 11203 4951 11209
rect 4893 11169 4905 11203
rect 4939 11200 4951 11203
rect 5074 11200 5080 11212
rect 4939 11172 5080 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 6454 11160 6460 11212
rect 6512 11200 6518 11212
rect 7466 11200 7472 11212
rect 6512 11172 7472 11200
rect 6512 11160 6518 11172
rect 7466 11160 7472 11172
rect 7524 11200 7530 11212
rect 9217 11203 9275 11209
rect 9217 11200 9229 11203
rect 7524 11172 9229 11200
rect 7524 11160 7530 11172
rect 9217 11169 9229 11172
rect 9263 11200 9275 11203
rect 9582 11200 9588 11212
rect 9263 11172 9588 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 9766 11160 9772 11212
rect 9824 11160 9830 11212
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3936 11104 3985 11132
rect 3936 11092 3942 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 4212 11104 4721 11132
rect 4212 11092 4218 11104
rect 4709 11101 4721 11104
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11132 5043 11135
rect 8110 11132 8116 11144
rect 5031 11104 8116 11132
rect 5031 11101 5043 11104
rect 4985 11095 5043 11101
rect 2590 10956 2596 11008
rect 2648 10996 2654 11008
rect 3510 10996 3516 11008
rect 2648 10968 3516 10996
rect 2648 10956 2654 10968
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 4246 10956 4252 11008
rect 4304 10956 4310 11008
rect 4341 10999 4399 11005
rect 4341 10965 4353 10999
rect 4387 10996 4399 10999
rect 4430 10996 4436 11008
rect 4387 10968 4436 10996
rect 4387 10965 4399 10968
rect 4341 10959 4399 10965
rect 4430 10956 4436 10968
rect 4488 10956 4494 11008
rect 4724 10996 4752 11095
rect 8110 11092 8116 11104
rect 8168 11132 8174 11144
rect 8662 11132 8668 11144
rect 8168 11104 8668 11132
rect 8168 11092 8174 11104
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 8754 11092 8760 11144
rect 8812 11132 8818 11144
rect 8938 11132 8944 11144
rect 8812 11104 8944 11132
rect 8812 11092 8818 11104
rect 8938 11092 8944 11104
rect 8996 11132 9002 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8996 11104 9137 11132
rect 8996 11092 9002 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 9784 11132 9812 11160
rect 9447 11104 9812 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 7282 11064 7288 11076
rect 6380 11036 7288 11064
rect 5994 10996 6000 11008
rect 4724 10968 6000 10996
rect 5994 10956 6000 10968
rect 6052 10996 6058 11008
rect 6380 10996 6408 11036
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 9324 11064 9352 11095
rect 8266 11036 9352 11064
rect 9585 11067 9643 11073
rect 6052 10968 6408 10996
rect 6052 10956 6058 10968
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 8110 10996 8116 11008
rect 6696 10968 8116 10996
rect 6696 10956 6702 10968
rect 8110 10956 8116 10968
rect 8168 10996 8174 11008
rect 8266 10996 8294 11036
rect 9585 11033 9597 11067
rect 9631 11064 9643 11067
rect 9766 11064 9772 11076
rect 9631 11036 9772 11064
rect 9631 11033 9643 11036
rect 9585 11027 9643 11033
rect 9766 11024 9772 11036
rect 9824 11064 9830 11076
rect 9876 11064 9904 11240
rect 9953 11237 9965 11271
rect 9999 11237 10011 11271
rect 9953 11231 10011 11237
rect 10045 11271 10103 11277
rect 10045 11237 10057 11271
rect 10091 11268 10103 11271
rect 10226 11268 10232 11280
rect 10091 11240 10232 11268
rect 10091 11237 10103 11240
rect 10045 11231 10103 11237
rect 9968 11200 9996 11231
rect 10226 11228 10232 11240
rect 10284 11228 10290 11280
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 12250 11268 12256 11280
rect 11756 11240 12256 11268
rect 11756 11228 11762 11240
rect 12250 11228 12256 11240
rect 12308 11228 12314 11280
rect 12360 11200 12388 11308
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 18509 11339 18567 11345
rect 18509 11336 18521 11339
rect 13596 11308 18521 11336
rect 13596 11296 13602 11308
rect 18509 11305 18521 11308
rect 18555 11305 18567 11339
rect 18509 11299 18567 11305
rect 15838 11228 15844 11280
rect 15896 11228 15902 11280
rect 14369 11203 14427 11209
rect 14369 11200 14381 11203
rect 9968 11172 11836 11200
rect 12360 11172 14381 11200
rect 10318 11092 10324 11144
rect 10376 11092 10382 11144
rect 11808 11132 11836 11172
rect 14369 11169 14381 11172
rect 14415 11169 14427 11203
rect 14369 11163 14427 11169
rect 16850 11160 16856 11212
rect 16908 11200 16914 11212
rect 18141 11203 18199 11209
rect 18141 11200 18153 11203
rect 16908 11172 18153 11200
rect 16908 11160 16914 11172
rect 18141 11169 18153 11172
rect 18187 11169 18199 11203
rect 18141 11163 18199 11169
rect 12526 11132 12532 11144
rect 11808 11104 12532 11132
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 14056 11104 14105 11132
rect 14056 11092 14062 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 17000 11104 18337 11132
rect 17000 11092 17006 11104
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 18325 11095 18383 11101
rect 9824 11036 9904 11064
rect 10597 11067 10655 11073
rect 9824 11024 9830 11036
rect 10597 11033 10609 11067
rect 10643 11033 10655 11067
rect 10597 11027 10655 11033
rect 8168 10968 8294 10996
rect 8168 10956 8174 10968
rect 9030 10956 9036 11008
rect 9088 10996 9094 11008
rect 10612 10996 10640 11027
rect 11054 11024 11060 11076
rect 11112 11024 11118 11076
rect 12250 11024 12256 11076
rect 12308 11064 12314 11076
rect 12345 11067 12403 11073
rect 12345 11064 12357 11067
rect 12308 11036 12357 11064
rect 12308 11024 12314 11036
rect 12345 11033 12357 11036
rect 12391 11033 12403 11067
rect 12345 11027 12403 11033
rect 14918 11024 14924 11076
rect 14976 11024 14982 11076
rect 9088 10968 10640 10996
rect 9088 10956 9094 10968
rect 11974 10956 11980 11008
rect 12032 10996 12038 11008
rect 14182 10996 14188 11008
rect 12032 10968 14188 10996
rect 12032 10956 12038 10968
rect 14182 10956 14188 10968
rect 14240 10956 14246 11008
rect 14550 10956 14556 11008
rect 14608 10996 14614 11008
rect 16390 10996 16396 11008
rect 14608 10968 16396 10996
rect 14608 10956 14614 10968
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 17310 10956 17316 11008
rect 17368 10996 17374 11008
rect 17494 10996 17500 11008
rect 17368 10968 17500 10996
rect 17368 10956 17374 10968
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 1104 10906 18860 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 17610 10906
rect 17662 10854 17674 10906
rect 17726 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 18860 10906
rect 1104 10832 18860 10854
rect 5442 10792 5448 10804
rect 2700 10764 5448 10792
rect 1670 10616 1676 10668
rect 1728 10656 1734 10668
rect 2700 10665 2728 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 7561 10795 7619 10801
rect 7561 10792 7573 10795
rect 5592 10764 7573 10792
rect 5592 10752 5598 10764
rect 7561 10761 7573 10764
rect 7607 10761 7619 10795
rect 11698 10792 11704 10804
rect 7561 10755 7619 10761
rect 9324 10764 11704 10792
rect 2777 10727 2835 10733
rect 2777 10693 2789 10727
rect 2823 10724 2835 10727
rect 5626 10724 5632 10736
rect 2823 10696 5632 10724
rect 2823 10693 2835 10696
rect 2777 10687 2835 10693
rect 5626 10684 5632 10696
rect 5684 10684 5690 10736
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 1728 10628 2697 10656
rect 1728 10616 1734 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 3602 10616 3608 10668
rect 3660 10616 3666 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5902 10656 5908 10668
rect 5592 10628 5908 10656
rect 5592 10616 5598 10628
rect 5902 10616 5908 10628
rect 5960 10656 5966 10668
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 5960 10628 7481 10656
rect 5960 10616 5966 10628
rect 7469 10625 7481 10628
rect 7515 10656 7527 10659
rect 8754 10656 8760 10668
rect 7515 10628 8760 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 9324 10588 9352 10764
rect 11698 10752 11704 10764
rect 11756 10792 11762 10804
rect 11974 10792 11980 10804
rect 11756 10764 11980 10792
rect 11756 10752 11762 10764
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 16206 10792 16212 10804
rect 14240 10764 16212 10792
rect 14240 10752 14246 10764
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 17678 10792 17684 10804
rect 17184 10764 17684 10792
rect 17184 10752 17190 10764
rect 17678 10752 17684 10764
rect 17736 10792 17742 10804
rect 17736 10764 18000 10792
rect 17736 10752 17742 10764
rect 9582 10684 9588 10736
rect 9640 10724 9646 10736
rect 16666 10724 16672 10736
rect 9640 10696 16672 10724
rect 9640 10684 9646 10696
rect 16666 10684 16672 10696
rect 16724 10724 16730 10736
rect 16850 10724 16856 10736
rect 16724 10696 16856 10724
rect 16724 10684 16730 10696
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 17218 10684 17224 10736
rect 17276 10684 17282 10736
rect 17405 10727 17463 10733
rect 17405 10693 17417 10727
rect 17451 10724 17463 10727
rect 17494 10724 17500 10736
rect 17451 10696 17500 10724
rect 17451 10693 17463 10696
rect 17405 10687 17463 10693
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 17972 10733 18000 10764
rect 17957 10727 18015 10733
rect 17957 10693 17969 10727
rect 18003 10693 18015 10727
rect 17957 10687 18015 10693
rect 18173 10727 18231 10733
rect 18173 10693 18185 10727
rect 18219 10724 18231 10727
rect 18690 10724 18696 10736
rect 18219 10696 18696 10724
rect 18219 10693 18231 10696
rect 18173 10687 18231 10693
rect 18690 10684 18696 10696
rect 18748 10684 18754 10736
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 17681 10659 17739 10665
rect 17681 10656 17693 10659
rect 10008 10628 17693 10656
rect 10008 10616 10014 10628
rect 17681 10625 17693 10628
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 2746 10560 9352 10588
rect 2406 10480 2412 10532
rect 2464 10520 2470 10532
rect 2746 10520 2774 10560
rect 9398 10548 9404 10600
rect 9456 10588 9462 10600
rect 14921 10591 14979 10597
rect 14921 10588 14933 10591
rect 9456 10560 14933 10588
rect 9456 10548 9462 10560
rect 14921 10557 14933 10560
rect 14967 10557 14979 10591
rect 14921 10551 14979 10557
rect 16666 10548 16672 10600
rect 16724 10588 16730 10600
rect 16942 10588 16948 10600
rect 16724 10560 16948 10588
rect 16724 10548 16730 10560
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 17586 10588 17592 10600
rect 17276 10560 17592 10588
rect 17276 10548 17282 10560
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 2464 10492 2774 10520
rect 2464 10480 2470 10492
rect 5258 10480 5264 10532
rect 5316 10520 5322 10532
rect 11054 10520 11060 10532
rect 5316 10492 11060 10520
rect 5316 10480 5322 10492
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 13170 10520 13176 10532
rect 11204 10492 13176 10520
rect 11204 10480 11210 10492
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 14182 10480 14188 10532
rect 14240 10520 14246 10532
rect 14458 10520 14464 10532
rect 14240 10492 14464 10520
rect 14240 10480 14246 10492
rect 14458 10480 14464 10492
rect 14516 10480 14522 10532
rect 15194 10480 15200 10532
rect 15252 10480 15258 10532
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 17494 10520 17500 10532
rect 15620 10492 17500 10520
rect 15620 10480 15626 10492
rect 17494 10480 17500 10492
rect 17552 10480 17558 10532
rect 18782 10520 18788 10532
rect 18156 10492 18788 10520
rect 18156 10464 18184 10492
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 3697 10455 3755 10461
rect 3697 10421 3709 10455
rect 3743 10452 3755 10455
rect 11514 10452 11520 10464
rect 3743 10424 11520 10452
rect 3743 10421 3755 10424
rect 3697 10415 3755 10421
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 15378 10412 15384 10464
rect 15436 10412 15442 10464
rect 16206 10412 16212 10464
rect 16264 10452 16270 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 16264 10424 17417 10452
rect 16264 10412 16270 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 18138 10412 18144 10464
rect 18196 10412 18202 10464
rect 18322 10412 18328 10464
rect 18380 10412 18386 10464
rect 1104 10362 18860 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 16950 10362
rect 17002 10310 17014 10362
rect 17066 10310 17078 10362
rect 17130 10310 17142 10362
rect 17194 10310 17206 10362
rect 17258 10310 18860 10362
rect 1104 10288 18860 10310
rect 6638 10248 6644 10260
rect 4540 10220 6644 10248
rect 4540 10121 4568 10220
rect 6638 10208 6644 10220
rect 6696 10248 6702 10260
rect 8294 10248 8300 10260
rect 6696 10220 8300 10248
rect 6696 10208 6702 10220
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 10870 10248 10876 10260
rect 9646 10220 10876 10248
rect 6914 10140 6920 10192
rect 6972 10180 6978 10192
rect 9646 10180 9674 10220
rect 10870 10208 10876 10220
rect 10928 10248 10934 10260
rect 15562 10248 15568 10260
rect 10928 10220 15568 10248
rect 10928 10208 10934 10220
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 15838 10248 15844 10260
rect 15703 10220 15844 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 6972 10152 9674 10180
rect 6972 10140 6978 10152
rect 13906 10140 13912 10192
rect 13964 10180 13970 10192
rect 13964 10152 16252 10180
rect 13964 10140 13970 10152
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 4614 10072 4620 10124
rect 4672 10072 4678 10124
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 4890 10112 4896 10124
rect 4847 10084 4896 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 5258 10072 5264 10124
rect 5316 10112 5322 10124
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 5316 10084 7389 10112
rect 5316 10072 5322 10084
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 7466 10072 7472 10124
rect 7524 10072 7530 10124
rect 7653 10115 7711 10121
rect 7653 10081 7665 10115
rect 7699 10112 7711 10115
rect 8202 10112 8208 10124
rect 7699 10084 8208 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 8202 10072 8208 10084
rect 8260 10112 8266 10124
rect 9582 10112 9588 10124
rect 8260 10084 9588 10112
rect 8260 10072 8266 10084
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 10597 10115 10655 10121
rect 10597 10112 10609 10115
rect 10468 10084 10609 10112
rect 10468 10072 10474 10084
rect 10597 10081 10609 10084
rect 10643 10112 10655 10115
rect 13998 10112 14004 10124
rect 10643 10084 14004 10112
rect 10643 10081 10655 10084
rect 10597 10075 10655 10081
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 16025 10115 16083 10121
rect 16025 10112 16037 10115
rect 14148 10084 16037 10112
rect 14148 10072 14154 10084
rect 16025 10081 16037 10084
rect 16071 10081 16083 10115
rect 16025 10075 16083 10081
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 4246 9936 4252 9988
rect 4304 9976 4310 9988
rect 4614 9976 4620 9988
rect 4304 9948 4620 9976
rect 4304 9936 4310 9948
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 4338 9868 4344 9920
rect 4396 9868 4402 9920
rect 4724 9908 4752 10007
rect 4982 10004 4988 10056
rect 5040 10004 5046 10056
rect 6730 10004 6736 10056
rect 6788 10004 6794 10056
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 7484 10044 7512 10072
rect 7064 10016 7512 10044
rect 7561 10047 7619 10053
rect 7064 10004 7070 10016
rect 7561 10013 7573 10047
rect 7607 10044 7619 10047
rect 8110 10044 8116 10056
rect 7607 10016 8116 10044
rect 7607 10013 7619 10016
rect 7561 10007 7619 10013
rect 5258 9936 5264 9988
rect 5316 9936 5322 9988
rect 5718 9936 5724 9988
rect 5776 9936 5782 9988
rect 6748 9976 6776 10004
rect 7576 9976 7604 10007
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 13872 10016 15853 10044
rect 13872 10004 13878 10016
rect 15841 10013 15853 10016
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 15930 10004 15936 10056
rect 15988 10004 15994 10056
rect 16114 10004 16120 10056
rect 16172 10004 16178 10056
rect 16224 10044 16252 10152
rect 16850 10140 16856 10192
rect 16908 10180 16914 10192
rect 17037 10183 17095 10189
rect 17037 10180 17049 10183
rect 16908 10152 17049 10180
rect 16908 10140 16914 10152
rect 17037 10149 17049 10152
rect 17083 10149 17095 10183
rect 17037 10143 17095 10149
rect 16942 10072 16948 10124
rect 17000 10112 17006 10124
rect 17586 10112 17592 10124
rect 17000 10084 17592 10112
rect 17000 10072 17006 10084
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 17313 10047 17371 10053
rect 17313 10044 17325 10047
rect 16224 10016 17325 10044
rect 17313 10013 17325 10016
rect 17359 10013 17371 10047
rect 17313 10007 17371 10013
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10044 17463 10047
rect 17678 10044 17684 10056
rect 17451 10016 17684 10044
rect 17451 10013 17463 10016
rect 17405 10007 17463 10013
rect 17678 10004 17684 10016
rect 17736 10044 17742 10056
rect 18046 10044 18052 10056
rect 17736 10016 18052 10044
rect 17736 10004 17742 10016
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 6748 9948 7604 9976
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 10594 9976 10600 9988
rect 8812 9948 10600 9976
rect 8812 9936 8818 9948
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 10873 9979 10931 9985
rect 10873 9945 10885 9979
rect 10919 9976 10931 9979
rect 11146 9976 11152 9988
rect 10919 9948 11152 9976
rect 10919 9945 10931 9948
rect 10873 9939 10931 9945
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 11256 9948 11362 9976
rect 5074 9908 5080 9920
rect 4724 9880 5080 9908
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 6546 9868 6552 9920
rect 6604 9908 6610 9920
rect 6733 9911 6791 9917
rect 6733 9908 6745 9911
rect 6604 9880 6745 9908
rect 6604 9868 6610 9880
rect 6733 9877 6745 9880
rect 6779 9877 6791 9911
rect 6733 9871 6791 9877
rect 7190 9868 7196 9920
rect 7248 9868 7254 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 8018 9908 8024 9920
rect 7524 9880 8024 9908
rect 7524 9868 7530 9880
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 11256 9908 11284 9948
rect 13722 9936 13728 9988
rect 13780 9976 13786 9988
rect 16132 9976 16160 10004
rect 13780 9948 16160 9976
rect 13780 9936 13786 9948
rect 16390 9936 16396 9988
rect 16448 9976 16454 9988
rect 16448 9948 17356 9976
rect 16448 9936 16454 9948
rect 9824 9880 11284 9908
rect 9824 9868 9830 9880
rect 12250 9868 12256 9920
rect 12308 9908 12314 9920
rect 12345 9911 12403 9917
rect 12345 9908 12357 9911
rect 12308 9880 12357 9908
rect 12308 9868 12314 9880
rect 12345 9877 12357 9880
rect 12391 9877 12403 9911
rect 12345 9871 12403 9877
rect 15838 9868 15844 9920
rect 15896 9908 15902 9920
rect 16206 9908 16212 9920
rect 15896 9880 16212 9908
rect 15896 9868 15902 9880
rect 16206 9868 16212 9880
rect 16264 9908 16270 9920
rect 17221 9911 17279 9917
rect 17221 9908 17233 9911
rect 16264 9880 17233 9908
rect 16264 9868 16270 9880
rect 17221 9877 17233 9880
rect 17267 9877 17279 9911
rect 17328 9908 17356 9948
rect 18138 9936 18144 9988
rect 18196 9936 18202 9988
rect 17589 9911 17647 9917
rect 17589 9908 17601 9911
rect 17328 9880 17601 9908
rect 17221 9871 17279 9877
rect 17589 9877 17601 9880
rect 17635 9877 17647 9911
rect 17589 9871 17647 9877
rect 18230 9868 18236 9920
rect 18288 9868 18294 9920
rect 1104 9818 18860 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 17610 9818
rect 17662 9766 17674 9818
rect 17726 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 18860 9818
rect 1104 9744 18860 9766
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 9030 9704 9036 9716
rect 3936 9676 8064 9704
rect 3936 9664 3942 9676
rect 1762 9596 1768 9648
rect 1820 9596 1826 9648
rect 6086 9596 6092 9648
rect 6144 9636 6150 9648
rect 8036 9636 8064 9676
rect 8266 9676 9036 9704
rect 8266 9636 8294 9676
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 10410 9704 10416 9716
rect 9232 9676 10416 9704
rect 9232 9636 9260 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 16390 9704 16396 9716
rect 16172 9676 16396 9704
rect 16172 9664 16178 9676
rect 16390 9664 16396 9676
rect 16448 9664 16454 9716
rect 10778 9636 10784 9648
rect 6144 9608 7222 9636
rect 8036 9608 8294 9636
rect 8588 9608 9260 9636
rect 10074 9608 10784 9636
rect 6144 9596 6150 9608
rect 1670 9528 1676 9580
rect 1728 9528 1734 9580
rect 5166 9528 5172 9580
rect 5224 9528 5230 9580
rect 8588 9577 8616 9608
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 14090 9636 14096 9648
rect 10888 9608 14096 9636
rect 8573 9571 8631 9577
rect 8573 9537 8585 9571
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 10888 9568 10916 9608
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 14277 9639 14335 9645
rect 14277 9605 14289 9639
rect 14323 9636 14335 9639
rect 14366 9636 14372 9648
rect 14323 9608 14372 9636
rect 14323 9605 14335 9608
rect 14277 9599 14335 9605
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 14458 9596 14464 9648
rect 14516 9636 14522 9648
rect 15654 9636 15660 9648
rect 14516 9608 15660 9636
rect 14516 9596 14522 9608
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 10284 9540 10916 9568
rect 10284 9528 10290 9540
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 11020 9540 12265 9568
rect 11020 9528 11026 9540
rect 12253 9537 12265 9540
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 5040 9472 6469 9500
rect 5040 9460 5046 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 7466 9500 7472 9512
rect 6779 9472 7472 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 5132 9336 5273 9364
rect 5132 9324 5138 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 6472 9364 6500 9463
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7742 9460 7748 9512
rect 7800 9500 7806 9512
rect 8205 9503 8263 9509
rect 8205 9500 8217 9503
rect 7800 9472 8217 9500
rect 7800 9460 7806 9472
rect 8205 9469 8217 9472
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 8846 9460 8852 9512
rect 8904 9460 8910 9512
rect 12268 9432 12296 9531
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 12492 9540 13461 9568
rect 12492 9528 12498 9540
rect 13449 9537 13461 9540
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 14826 9568 14832 9580
rect 14608 9540 14832 9568
rect 14608 9528 14614 9540
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12400 9472 14320 9500
rect 12400 9460 12406 9472
rect 14292 9441 14320 9472
rect 14277 9435 14335 9441
rect 12268 9404 14228 9432
rect 8294 9364 8300 9376
rect 6472 9336 8300 9364
rect 5261 9327 5319 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 9858 9324 9864 9376
rect 9916 9364 9922 9376
rect 10321 9367 10379 9373
rect 10321 9364 10333 9367
rect 9916 9336 10333 9364
rect 9916 9324 9922 9336
rect 10321 9333 10333 9336
rect 10367 9364 10379 9367
rect 10870 9364 10876 9376
rect 10367 9336 10876 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 12345 9367 12403 9373
rect 12345 9364 12357 9367
rect 11296 9336 12357 9364
rect 11296 9324 11302 9336
rect 12345 9333 12357 9336
rect 12391 9333 12403 9367
rect 12345 9327 12403 9333
rect 13633 9367 13691 9373
rect 13633 9333 13645 9367
rect 13679 9364 13691 9367
rect 13814 9364 13820 9376
rect 13679 9336 13820 9364
rect 13679 9333 13691 9336
rect 13633 9327 13691 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 14200 9364 14228 9404
rect 14277 9401 14289 9435
rect 14323 9401 14335 9435
rect 14277 9395 14335 9401
rect 15470 9364 15476 9376
rect 14200 9336 15476 9364
rect 15470 9324 15476 9336
rect 15528 9364 15534 9376
rect 15838 9364 15844 9376
rect 15528 9336 15844 9364
rect 15528 9324 15534 9336
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 1104 9274 18860 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 16950 9274
rect 17002 9222 17014 9274
rect 17066 9222 17078 9274
rect 17130 9222 17142 9274
rect 17194 9222 17206 9274
rect 17258 9222 18860 9274
rect 1104 9200 18860 9222
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 3476 9132 7052 9160
rect 3476 9120 3482 9132
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 6917 9095 6975 9101
rect 6917 9092 6929 9095
rect 3568 9064 6929 9092
rect 3568 9052 3574 9064
rect 6917 9061 6929 9064
rect 6963 9061 6975 9095
rect 7024 9092 7052 9132
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 13909 9163 13967 9169
rect 13909 9160 13921 9163
rect 7432 9132 13921 9160
rect 7432 9120 7438 9132
rect 13909 9129 13921 9132
rect 13955 9129 13967 9163
rect 13909 9123 13967 9129
rect 7653 9095 7711 9101
rect 7653 9092 7665 9095
rect 7024 9064 7665 9092
rect 6917 9055 6975 9061
rect 7653 9061 7665 9064
rect 7699 9061 7711 9095
rect 7653 9055 7711 9061
rect 7834 9052 7840 9104
rect 7892 9092 7898 9104
rect 7892 9064 8248 9092
rect 7892 9052 7898 9064
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 6454 9024 6460 9036
rect 5132 8996 6460 9024
rect 5132 8984 5138 8996
rect 6454 8984 6460 8996
rect 6512 9024 6518 9036
rect 6758 9027 6816 9033
rect 6758 9024 6770 9027
rect 6512 8996 6770 9024
rect 6512 8984 6518 8996
rect 6758 8993 6770 8996
rect 6804 8993 6816 9027
rect 6758 8987 6816 8993
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7852 9024 7880 9052
rect 7064 8996 7880 9024
rect 7064 8984 7070 8996
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 8220 9033 8248 9064
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 9582 9092 9588 9104
rect 8444 9064 9588 9092
rect 8444 9052 8450 9064
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 11054 9052 11060 9104
rect 11112 9092 11118 9104
rect 11514 9092 11520 9104
rect 11112 9064 11520 9092
rect 11112 9052 11118 9064
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 8113 9027 8171 9033
rect 8113 9024 8125 9027
rect 7984 8996 8125 9024
rect 7984 8984 7990 8996
rect 8113 8993 8125 8996
rect 8159 8993 8171 9027
rect 8113 8987 8171 8993
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 8993 8263 9027
rect 13722 9024 13728 9036
rect 8205 8987 8263 8993
rect 8312 8996 13728 9024
rect 1489 8959 1547 8965
rect 1489 8925 1501 8959
rect 1535 8956 1547 8959
rect 2958 8956 2964 8968
rect 1535 8928 2964 8956
rect 1535 8925 1547 8928
rect 1489 8919 1547 8925
rect 2958 8916 2964 8928
rect 3016 8956 3022 8968
rect 3970 8956 3976 8968
rect 3016 8928 3976 8956
rect 3016 8916 3022 8928
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 6380 8928 6653 8956
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 6086 8888 6092 8900
rect 5040 8860 6092 8888
rect 5040 8848 5046 8860
rect 6086 8848 6092 8860
rect 6144 8888 6150 8900
rect 6380 8888 6408 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 7282 8916 7288 8968
rect 7340 8956 7346 8968
rect 8312 8956 8340 8996
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 7340 8928 8340 8956
rect 7340 8916 7346 8928
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8720 8928 8953 8956
rect 8720 8916 8726 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9582 8956 9588 8968
rect 9263 8928 9588 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 11848 8928 12173 8956
rect 11848 8916 11854 8928
rect 12161 8925 12173 8928
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 14921 8959 14979 8965
rect 14921 8925 14933 8959
rect 14967 8956 14979 8959
rect 18230 8956 18236 8968
rect 14967 8928 18236 8956
rect 14967 8925 14979 8928
rect 14921 8919 14979 8925
rect 6144 8860 6408 8888
rect 8021 8891 8079 8897
rect 6144 8848 6150 8860
rect 8021 8857 8033 8891
rect 8067 8888 8079 8891
rect 8754 8888 8760 8900
rect 8067 8860 8760 8888
rect 8067 8857 8079 8860
rect 8021 8851 8079 8857
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9306 8888 9312 8900
rect 9088 8860 9312 8888
rect 9088 8848 9094 8860
rect 9306 8848 9312 8860
rect 9364 8848 9370 8900
rect 11054 8848 11060 8900
rect 11112 8888 11118 8900
rect 12437 8891 12495 8897
rect 12437 8888 12449 8891
rect 11112 8860 12449 8888
rect 11112 8848 11118 8860
rect 12437 8857 12449 8860
rect 12483 8857 12495 8891
rect 12437 8851 12495 8857
rect 13078 8848 13084 8900
rect 13136 8848 13142 8900
rect 934 8780 940 8832
rect 992 8820 998 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 992 8792 1593 8820
rect 992 8780 998 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 6549 8823 6607 8829
rect 6549 8789 6561 8823
rect 6595 8820 6607 8823
rect 8386 8820 8392 8832
rect 6595 8792 8392 8820
rect 6595 8789 6607 8792
rect 6549 8783 6607 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 8536 8792 9137 8820
rect 8536 8780 8542 8792
rect 9125 8789 9137 8792
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 9398 8780 9404 8832
rect 9456 8820 9462 8832
rect 9493 8823 9551 8829
rect 9493 8820 9505 8823
rect 9456 8792 9505 8820
rect 9456 8780 9462 8792
rect 9493 8789 9505 8792
rect 9539 8789 9551 8823
rect 9493 8783 9551 8789
rect 10318 8780 10324 8832
rect 10376 8820 10382 8832
rect 12526 8820 12532 8832
rect 10376 8792 12532 8820
rect 10376 8780 10382 8792
rect 12526 8780 12532 8792
rect 12584 8820 12590 8832
rect 14936 8820 14964 8919
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 15749 8891 15807 8897
rect 15749 8857 15761 8891
rect 15795 8888 15807 8891
rect 15838 8888 15844 8900
rect 15795 8860 15844 8888
rect 15795 8857 15807 8860
rect 15749 8851 15807 8857
rect 15838 8848 15844 8860
rect 15896 8848 15902 8900
rect 12584 8792 14964 8820
rect 12584 8780 12590 8792
rect 1104 8730 18860 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 17610 8730
rect 17662 8678 17674 8730
rect 17726 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 18860 8730
rect 1104 8656 18860 8678
rect 3786 8576 3792 8628
rect 3844 8576 3850 8628
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 5500 8588 10609 8616
rect 5500 8576 5506 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 10597 8579 10655 8585
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 13725 8619 13783 8625
rect 13725 8616 13737 8619
rect 11204 8588 13737 8616
rect 11204 8576 11210 8588
rect 13725 8585 13737 8588
rect 13771 8585 13783 8619
rect 13725 8579 13783 8585
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 8570 8548 8576 8560
rect 8260 8520 8576 8548
rect 8260 8508 8266 8520
rect 8570 8508 8576 8520
rect 8628 8548 8634 8560
rect 8628 8520 10640 8548
rect 8628 8508 8634 8520
rect 3234 8440 3240 8492
rect 3292 8480 3298 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3292 8452 3433 8480
rect 3292 8440 3298 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 3970 8480 3976 8492
rect 3651 8452 3976 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 10612 8480 10640 8520
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 13998 8548 14004 8560
rect 11572 8520 14004 8548
rect 11572 8508 11578 8520
rect 13998 8508 14004 8520
rect 14056 8548 14062 8560
rect 15930 8548 15936 8560
rect 14056 8520 15936 8548
rect 14056 8508 14062 8520
rect 15930 8508 15936 8520
rect 15988 8508 15994 8560
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 10612 8452 17693 8480
rect 17681 8449 17693 8452
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 6454 8412 6460 8424
rect 4948 8384 6460 8412
rect 4948 8372 4954 8384
rect 6454 8372 6460 8384
rect 6512 8412 6518 8424
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 6512 8384 6561 8412
rect 6512 8372 6518 8384
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 7006 8372 7012 8424
rect 7064 8372 7070 8424
rect 7374 8412 7380 8424
rect 7432 8421 7438 8424
rect 7432 8415 7460 8421
rect 7116 8384 7380 8412
rect 5902 8304 5908 8356
rect 5960 8344 5966 8356
rect 7024 8344 7052 8372
rect 5960 8316 7052 8344
rect 5960 8304 5966 8316
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 7116 8276 7144 8384
rect 7374 8372 7380 8384
rect 7448 8381 7460 8415
rect 7432 8375 7460 8381
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 7607 8384 7972 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 7432 8372 7438 8375
rect 6144 8248 7144 8276
rect 7944 8276 7972 8384
rect 8110 8372 8116 8424
rect 8168 8412 8174 8424
rect 8168 8384 12388 8412
rect 8168 8372 8174 8384
rect 12360 8356 12388 8384
rect 13814 8372 13820 8424
rect 13872 8412 13878 8424
rect 13909 8415 13967 8421
rect 13909 8412 13921 8415
rect 13872 8384 13921 8412
rect 13872 8372 13878 8384
rect 13909 8381 13921 8384
rect 13955 8381 13967 8415
rect 13909 8375 13967 8381
rect 13998 8372 14004 8424
rect 14056 8372 14062 8424
rect 14090 8372 14096 8424
rect 14148 8372 14154 8424
rect 14185 8415 14243 8421
rect 14185 8381 14197 8415
rect 14231 8381 14243 8415
rect 14185 8375 14243 8381
rect 8202 8304 8208 8356
rect 8260 8304 8266 8356
rect 10520 8316 10732 8344
rect 8386 8276 8392 8288
rect 7944 8248 8392 8276
rect 6144 8236 6150 8248
rect 8386 8236 8392 8248
rect 8444 8276 8450 8288
rect 8754 8276 8760 8288
rect 8444 8248 8760 8276
rect 8444 8236 8450 8248
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 10520 8276 10548 8316
rect 8904 8248 10548 8276
rect 10704 8276 10732 8316
rect 12342 8304 12348 8356
rect 12400 8344 12406 8356
rect 14200 8344 14228 8375
rect 12400 8316 14228 8344
rect 12400 8304 12406 8316
rect 15102 8304 15108 8356
rect 15160 8344 15166 8356
rect 17957 8347 18015 8353
rect 17957 8344 17969 8347
rect 15160 8316 17969 8344
rect 15160 8304 15166 8316
rect 17957 8313 17969 8316
rect 18003 8313 18015 8347
rect 17957 8307 18015 8313
rect 18138 8304 18144 8356
rect 18196 8304 18202 8356
rect 14826 8276 14832 8288
rect 10704 8248 14832 8276
rect 8904 8236 8910 8248
rect 14826 8236 14832 8248
rect 14884 8236 14890 8288
rect 1104 8186 18860 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 16950 8186
rect 17002 8134 17014 8186
rect 17066 8134 17078 8186
rect 17130 8134 17142 8186
rect 17194 8134 17206 8186
rect 17258 8134 18860 8186
rect 1104 8112 18860 8134
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 6273 8075 6331 8081
rect 6273 8072 6285 8075
rect 5316 8044 6285 8072
rect 5316 8032 5322 8044
rect 6273 8041 6285 8044
rect 6319 8041 6331 8075
rect 6273 8035 6331 8041
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 7006 8072 7012 8084
rect 6788 8044 7012 8072
rect 6788 8032 6794 8044
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 11057 8075 11115 8081
rect 11057 8041 11069 8075
rect 11103 8072 11115 8075
rect 15286 8072 15292 8084
rect 11103 8044 15292 8072
rect 11103 8041 11115 8044
rect 11057 8035 11115 8041
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 2869 8007 2927 8013
rect 2869 7973 2881 8007
rect 2915 8004 2927 8007
rect 9766 8004 9772 8016
rect 2915 7976 9772 8004
rect 2915 7973 2927 7976
rect 2869 7967 2927 7973
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 10137 8007 10195 8013
rect 10137 7973 10149 8007
rect 10183 8004 10195 8007
rect 16298 8004 16304 8016
rect 10183 7976 16304 8004
rect 10183 7973 10195 7976
rect 10137 7967 10195 7973
rect 16298 7964 16304 7976
rect 16356 7964 16362 8016
rect 6580 7908 6914 7936
rect 6580 7880 6608 7908
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 6546 7878 6552 7880
rect 6472 7877 6552 7878
rect 2777 7871 2835 7877
rect 2777 7868 2789 7871
rect 2464 7840 2789 7868
rect 2464 7828 2470 7840
rect 2777 7837 2789 7840
rect 2823 7837 2835 7871
rect 2777 7831 2835 7837
rect 6457 7871 6552 7877
rect 6457 7837 6469 7871
rect 6503 7850 6552 7871
rect 6503 7837 6515 7850
rect 6457 7831 6515 7837
rect 6546 7828 6552 7850
rect 6604 7828 6610 7880
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 6886 7868 6914 7908
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 8812 7908 10241 7936
rect 8812 7896 8818 7908
rect 10229 7905 10241 7908
rect 10275 7905 10287 7939
rect 12434 7936 12440 7948
rect 10229 7899 10287 7905
rect 10336 7908 12440 7936
rect 10336 7868 10364 7908
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 6886 7840 10364 7868
rect 10962 7828 10968 7880
rect 11020 7828 11026 7880
rect 9766 7760 9772 7812
rect 9824 7800 9830 7812
rect 17310 7800 17316 7812
rect 9824 7772 17316 7800
rect 9824 7760 9830 7772
rect 17310 7760 17316 7772
rect 17368 7760 17374 7812
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 6641 7735 6699 7741
rect 6641 7732 6653 7735
rect 5592 7704 6653 7732
rect 5592 7692 5598 7704
rect 6641 7701 6653 7704
rect 6687 7701 6699 7735
rect 6641 7695 6699 7701
rect 1104 7642 18860 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 17610 7642
rect 17662 7590 17674 7642
rect 17726 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 18860 7642
rect 1104 7568 18860 7590
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 11977 7531 12035 7537
rect 11977 7528 11989 7531
rect 3200 7500 11989 7528
rect 3200 7488 3206 7500
rect 11977 7497 11989 7500
rect 12023 7497 12035 7531
rect 11977 7491 12035 7497
rect 7374 7460 7380 7472
rect 6288 7432 7380 7460
rect 6288 7426 6316 7432
rect 5350 7352 5356 7404
rect 5408 7392 5414 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 5408 7364 5457 7392
rect 5408 7352 5414 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 5718 7392 5724 7404
rect 5445 7355 5503 7361
rect 5552 7364 5724 7392
rect 5552 7333 5580 7364
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 5810 7352 5816 7404
rect 5868 7392 5874 7404
rect 6196 7401 6316 7426
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 15010 7460 15016 7472
rect 9508 7432 15016 7460
rect 5905 7395 5963 7401
rect 5905 7392 5917 7395
rect 5868 7364 5917 7392
rect 5868 7352 5874 7364
rect 5905 7361 5917 7364
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 6089 7395 6147 7401
rect 6089 7361 6101 7395
rect 6135 7361 6147 7395
rect 6089 7355 6147 7361
rect 6181 7398 6316 7401
rect 6181 7395 6239 7398
rect 6181 7361 6193 7395
rect 6227 7361 6239 7395
rect 6181 7355 6239 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 6914 7392 6920 7404
rect 6871 7364 6920 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 5537 7327 5595 7333
rect 5537 7293 5549 7327
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 5644 7296 6040 7324
rect 3970 7216 3976 7268
rect 4028 7256 4034 7268
rect 5644 7256 5672 7296
rect 4028 7228 5672 7256
rect 4028 7216 4034 7228
rect 5718 7216 5724 7268
rect 5776 7256 5782 7268
rect 5813 7259 5871 7265
rect 5813 7256 5825 7259
rect 5776 7228 5825 7256
rect 5776 7216 5782 7228
rect 5813 7225 5825 7228
rect 5859 7225 5871 7259
rect 5813 7219 5871 7225
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 4580 7160 5917 7188
rect 4580 7148 4586 7160
rect 5905 7157 5917 7160
rect 5951 7157 5963 7191
rect 6012 7188 6040 7296
rect 6104 7256 6132 7355
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7392 7711 7395
rect 8018 7392 8024 7404
rect 7699 7364 8024 7392
rect 7699 7361 7711 7364
rect 7653 7355 7711 7361
rect 8018 7352 8024 7364
rect 8076 7392 8082 7404
rect 9508 7392 9536 7432
rect 15010 7420 15016 7432
rect 15068 7420 15074 7472
rect 8076 7364 9536 7392
rect 8076 7352 8082 7364
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 11204 7364 12173 7392
rect 11204 7352 11210 7364
rect 12161 7361 12173 7364
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 12434 7352 12440 7404
rect 12492 7352 12498 7404
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 17402 7392 17408 7404
rect 13504 7364 17408 7392
rect 13504 7352 13510 7364
rect 17402 7352 17408 7364
rect 17460 7392 17466 7404
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 17460 7364 17877 7392
rect 17460 7352 17466 7364
rect 17865 7361 17877 7364
rect 17911 7361 17923 7395
rect 17865 7355 17923 7361
rect 6546 7284 6552 7336
rect 6604 7284 6610 7336
rect 6638 7284 6644 7336
rect 6696 7284 6702 7336
rect 6730 7284 6736 7336
rect 6788 7284 6794 7336
rect 12345 7327 12403 7333
rect 12345 7293 12357 7327
rect 12391 7324 12403 7327
rect 16850 7324 16856 7336
rect 12391 7296 16856 7324
rect 12391 7293 12403 7296
rect 12345 7287 12403 7293
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 7006 7256 7012 7268
rect 6104 7228 7012 7256
rect 7006 7216 7012 7228
rect 7064 7216 7070 7268
rect 7098 7216 7104 7268
rect 7156 7256 7162 7268
rect 12986 7256 12992 7268
rect 7156 7228 12992 7256
rect 7156 7216 7162 7228
rect 12986 7216 12992 7228
rect 13044 7216 13050 7268
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 6012 7160 6377 7188
rect 5905 7151 5963 7157
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 7024 7188 7052 7216
rect 7558 7188 7564 7200
rect 7024 7160 7564 7188
rect 6365 7151 6423 7157
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 7837 7191 7895 7197
rect 7837 7157 7849 7191
rect 7883 7188 7895 7191
rect 8018 7188 8024 7200
rect 7883 7160 8024 7188
rect 7883 7157 7895 7160
rect 7837 7151 7895 7157
rect 8018 7148 8024 7160
rect 8076 7188 8082 7200
rect 8294 7188 8300 7200
rect 8076 7160 8300 7188
rect 8076 7148 8082 7160
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 16574 7188 16580 7200
rect 10928 7160 16580 7188
rect 10928 7148 10934 7160
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 17310 7148 17316 7200
rect 17368 7188 17374 7200
rect 17957 7191 18015 7197
rect 17957 7188 17969 7191
rect 17368 7160 17969 7188
rect 17368 7148 17374 7160
rect 17957 7157 17969 7160
rect 18003 7157 18015 7191
rect 17957 7151 18015 7157
rect 1104 7098 18860 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 16950 7098
rect 17002 7046 17014 7098
rect 17066 7046 17078 7098
rect 17130 7046 17142 7098
rect 17194 7046 17206 7098
rect 17258 7046 18860 7098
rect 1104 7024 18860 7046
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 5810 6984 5816 6996
rect 3384 6956 5816 6984
rect 3384 6944 3390 6956
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 10042 6984 10048 6996
rect 5920 6956 10048 6984
rect 5350 6876 5356 6928
rect 5408 6916 5414 6928
rect 5920 6916 5948 6956
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 11422 6944 11428 6996
rect 11480 6984 11486 6996
rect 11882 6984 11888 6996
rect 11480 6956 11888 6984
rect 11480 6944 11486 6956
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 13722 6984 13728 6996
rect 12400 6956 13728 6984
rect 12400 6944 12406 6956
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 5408 6888 5948 6916
rect 5408 6876 5414 6888
rect 5994 6876 6000 6928
rect 6052 6916 6058 6928
rect 8754 6916 8760 6928
rect 6052 6888 8760 6916
rect 6052 6876 6058 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 12434 6876 12440 6928
rect 12492 6916 12498 6928
rect 13446 6916 13452 6928
rect 12492 6888 13452 6916
rect 12492 6876 12498 6888
rect 13446 6876 13452 6888
rect 13504 6876 13510 6928
rect 3602 6808 3608 6860
rect 3660 6848 3666 6860
rect 4246 6848 4252 6860
rect 3660 6820 4252 6848
rect 3660 6808 3666 6820
rect 4246 6808 4252 6820
rect 4304 6848 4310 6860
rect 4304 6820 5948 6848
rect 4304 6808 4310 6820
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 5810 6780 5816 6792
rect 4672 6752 5816 6780
rect 4672 6740 4678 6752
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 5920 6780 5948 6820
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 12986 6848 12992 6860
rect 7616 6820 12992 6848
rect 7616 6808 7622 6820
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 16448 6820 17417 6848
rect 16448 6808 16454 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17405 6811 17463 6817
rect 10410 6780 10416 6792
rect 5920 6752 10416 6780
rect 10410 6740 10416 6752
rect 10468 6780 10474 6792
rect 12342 6780 12348 6792
rect 10468 6752 12348 6780
rect 10468 6740 10474 6752
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 15896 6752 17325 6780
rect 15896 6740 15902 6752
rect 17313 6749 17325 6752
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6780 18015 6783
rect 18003 6752 18184 6780
rect 18003 6749 18015 6752
rect 17957 6743 18015 6749
rect 3786 6672 3792 6724
rect 3844 6712 3850 6724
rect 6730 6712 6736 6724
rect 3844 6684 6736 6712
rect 3844 6672 3850 6684
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 14274 6712 14280 6724
rect 8720 6684 14280 6712
rect 8720 6672 8726 6684
rect 14274 6672 14280 6684
rect 14332 6712 14338 6724
rect 14642 6712 14648 6724
rect 14332 6684 14648 6712
rect 14332 6672 14338 6684
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 18049 6715 18107 6721
rect 18049 6712 18061 6715
rect 16816 6684 18061 6712
rect 16816 6672 16822 6684
rect 18049 6681 18061 6684
rect 18095 6681 18107 6715
rect 18049 6675 18107 6681
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 7650 6644 7656 6656
rect 5868 6616 7656 6644
rect 5868 6604 5874 6616
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 13630 6604 13636 6656
rect 13688 6644 13694 6656
rect 18156 6644 18184 6752
rect 13688 6616 18184 6644
rect 13688 6604 13694 6616
rect 1104 6554 18860 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 17610 6554
rect 17662 6502 17674 6554
rect 17726 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 18860 6554
rect 1104 6480 18860 6502
rect 6086 6440 6092 6452
rect 3252 6412 6092 6440
rect 2406 6372 2412 6384
rect 1964 6344 2412 6372
rect 1964 6316 1992 6344
rect 2406 6332 2412 6344
rect 2464 6332 2470 6384
rect 2866 6332 2872 6384
rect 2924 6372 2930 6384
rect 3050 6372 3056 6384
rect 2924 6344 3056 6372
rect 2924 6332 2930 6344
rect 3050 6332 3056 6344
rect 3108 6332 3114 6384
rect 1486 6264 1492 6316
rect 1544 6264 1550 6316
rect 1946 6264 1952 6316
rect 2004 6264 2010 6316
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6304 3019 6307
rect 3142 6304 3148 6316
rect 3007 6276 3148 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 2406 6236 2412 6248
rect 2363 6208 2412 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2041 6171 2099 6177
rect 2041 6137 2053 6171
rect 2087 6168 2099 6171
rect 2516 6168 2544 6267
rect 2792 6236 2820 6267
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3252 6313 3280 6412
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6178 6400 6184 6452
rect 6236 6400 6242 6452
rect 8018 6400 8024 6452
rect 8076 6400 8082 6452
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 14001 6443 14059 6449
rect 14001 6440 14013 6443
rect 10744 6412 14013 6440
rect 10744 6400 10750 6412
rect 14001 6409 14013 6412
rect 14047 6409 14059 6443
rect 14001 6403 14059 6409
rect 3421 6375 3479 6381
rect 3421 6341 3433 6375
rect 3467 6372 3479 6375
rect 3602 6372 3608 6384
rect 3467 6344 3608 6372
rect 3467 6341 3479 6344
rect 3421 6335 3479 6341
rect 3602 6332 3608 6344
rect 3660 6332 3666 6384
rect 4614 6372 4620 6384
rect 3896 6344 4620 6372
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6273 3295 6307
rect 3237 6267 3295 6273
rect 3510 6264 3516 6316
rect 3568 6264 3574 6316
rect 3602 6236 3608 6248
rect 2792 6208 3608 6236
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3053 6171 3111 6177
rect 2087 6140 2452 6168
rect 2516 6140 3004 6168
rect 2087 6137 2099 6140
rect 2041 6131 2099 6137
rect 934 6060 940 6112
rect 992 6100 998 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 992 6072 1593 6100
rect 992 6060 998 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 2424 6100 2452 6140
rect 2866 6100 2872 6112
rect 2424 6072 2872 6100
rect 1581 6063 1639 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 2976 6100 3004 6140
rect 3053 6137 3065 6171
rect 3099 6168 3111 6171
rect 3896 6168 3924 6344
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 4706 6332 4712 6384
rect 4764 6332 4770 6384
rect 6822 6372 6828 6384
rect 5934 6344 6828 6372
rect 6822 6332 6828 6344
rect 6880 6332 6886 6384
rect 8036 6372 8064 6400
rect 11606 6372 11612 6384
rect 7576 6344 8064 6372
rect 9062 6344 11612 6372
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 3988 6236 4016 6267
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4433 6307 4491 6313
rect 4433 6304 4445 6307
rect 4304 6276 4445 6304
rect 4304 6264 4310 6276
rect 4433 6273 4445 6276
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 5994 6264 6000 6316
rect 6052 6264 6058 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 7576 6313 7604 6344
rect 11606 6332 11612 6344
rect 11664 6332 11670 6384
rect 15194 6372 15200 6384
rect 12406 6344 15200 6372
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6236 6276 6561 6304
rect 6236 6264 6242 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 6549 6267 6607 6273
rect 6748 6276 7573 6304
rect 6012 6236 6040 6264
rect 3988 6208 6040 6236
rect 6638 6196 6644 6248
rect 6696 6196 6702 6248
rect 3099 6140 3924 6168
rect 3099 6137 3111 6140
rect 3053 6131 3111 6137
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 6748 6168 6776 6276
rect 7561 6273 7573 6276
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 12406 6304 12434 6344
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 9180 6276 12434 6304
rect 13725 6307 13783 6313
rect 9180 6264 9186 6276
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 14458 6304 14464 6316
rect 13771 6276 14464 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 18104 6276 18245 6304
rect 18104 6264 18110 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 10134 6236 10140 6248
rect 7883 6208 10140 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 13078 6236 13084 6248
rect 10652 6208 13084 6236
rect 10652 6196 10658 6208
rect 13078 6196 13084 6208
rect 13136 6236 13142 6248
rect 13630 6236 13636 6248
rect 13136 6208 13636 6236
rect 13136 6196 13142 6208
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 14001 6239 14059 6245
rect 14001 6205 14013 6239
rect 14047 6236 14059 6239
rect 16022 6236 16028 6248
rect 14047 6208 16028 6236
rect 14047 6205 14059 6208
rect 14001 6199 14059 6205
rect 6052 6140 6776 6168
rect 6840 6140 7696 6168
rect 6052 6128 6058 6140
rect 3786 6100 3792 6112
rect 2976 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6100 4215 6103
rect 6840 6100 6868 6140
rect 4203 6072 6868 6100
rect 6917 6103 6975 6109
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 6917 6069 6929 6103
rect 6963 6100 6975 6103
rect 7466 6100 7472 6112
rect 6963 6072 7472 6100
rect 6963 6069 6975 6072
rect 6917 6063 6975 6069
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7668 6100 7696 6140
rect 11882 6128 11888 6180
rect 11940 6168 11946 6180
rect 12618 6168 12624 6180
rect 11940 6140 12624 6168
rect 11940 6128 11946 6140
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 14016 6168 14044 6199
rect 16022 6196 16028 6208
rect 16080 6196 16086 6248
rect 13648 6140 14044 6168
rect 13648 6112 13676 6140
rect 18414 6128 18420 6180
rect 18472 6128 18478 6180
rect 8294 6100 8300 6112
rect 7668 6072 8300 6100
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 9306 6060 9312 6112
rect 9364 6060 9370 6112
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 11514 6100 11520 6112
rect 9456 6072 11520 6100
rect 9456 6060 9462 6072
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 13630 6060 13636 6112
rect 13688 6060 13694 6112
rect 13817 6103 13875 6109
rect 13817 6069 13829 6103
rect 13863 6100 13875 6103
rect 14550 6100 14556 6112
rect 13863 6072 14556 6100
rect 13863 6069 13875 6072
rect 13817 6063 13875 6069
rect 14550 6060 14556 6072
rect 14608 6100 14614 6112
rect 15102 6100 15108 6112
rect 14608 6072 15108 6100
rect 14608 6060 14614 6072
rect 15102 6060 15108 6072
rect 15160 6060 15166 6112
rect 1104 6010 18860 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 16950 6010
rect 17002 5958 17014 6010
rect 17066 5958 17078 6010
rect 17130 5958 17142 6010
rect 17194 5958 17206 6010
rect 17258 5958 18860 6010
rect 1104 5936 18860 5958
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 3973 5899 4031 5905
rect 3973 5896 3985 5899
rect 3936 5868 3985 5896
rect 3936 5856 3942 5868
rect 3973 5865 3985 5868
rect 4019 5865 4031 5899
rect 7282 5896 7288 5908
rect 3973 5859 4031 5865
rect 5276 5868 7288 5896
rect 3602 5788 3608 5840
rect 3660 5828 3666 5840
rect 3660 5800 4660 5828
rect 3660 5788 3666 5800
rect 4522 5760 4528 5772
rect 3988 5732 4528 5760
rect 3988 5701 4016 5732
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 4632 5692 4660 5800
rect 5276 5692 5304 5868
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7377 5899 7435 5905
rect 7377 5865 7389 5899
rect 7423 5896 7435 5899
rect 9122 5896 9128 5908
rect 7423 5868 9128 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 11388 5868 15669 5896
rect 11388 5856 11394 5868
rect 15657 5865 15669 5868
rect 15703 5865 15715 5899
rect 15657 5859 15715 5865
rect 8018 5828 8024 5840
rect 7484 5800 8024 5828
rect 5718 5720 5724 5772
rect 5776 5720 5782 5772
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 7484 5760 7512 5800
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 9398 5828 9404 5840
rect 8168 5800 9404 5828
rect 8168 5788 8174 5800
rect 9398 5788 9404 5800
rect 9456 5788 9462 5840
rect 14918 5828 14924 5840
rect 9968 5800 14924 5828
rect 6236 5732 7512 5760
rect 7561 5763 7619 5769
rect 6236 5720 6242 5732
rect 7561 5729 7573 5763
rect 7607 5760 7619 5763
rect 9030 5760 9036 5772
rect 7607 5732 8064 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 4203 5664 5304 5692
rect 5445 5695 5503 5701
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 5445 5661 5457 5695
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 2746 5596 4200 5624
rect 1486 5516 1492 5568
rect 1544 5556 1550 5568
rect 2746 5556 2774 5596
rect 1544 5528 2774 5556
rect 4172 5556 4200 5596
rect 4246 5584 4252 5636
rect 4304 5624 4310 5636
rect 5460 5624 5488 5655
rect 6822 5652 6828 5704
rect 6880 5652 6886 5704
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7432 5664 7665 5692
rect 7432 5652 7438 5664
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 5994 5624 6000 5636
rect 4304 5596 6000 5624
rect 4304 5584 4310 5596
rect 5994 5584 6000 5596
rect 6052 5584 6058 5636
rect 7282 5624 7288 5636
rect 7116 5596 7288 5624
rect 7116 5556 7144 5596
rect 7282 5584 7288 5596
rect 7340 5584 7346 5636
rect 7558 5584 7564 5636
rect 7616 5624 7622 5636
rect 7760 5624 7788 5655
rect 7834 5652 7840 5704
rect 7892 5652 7898 5704
rect 8036 5692 8064 5732
rect 8220 5732 9036 5760
rect 8220 5692 8248 5732
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 9674 5720 9680 5772
rect 9732 5720 9738 5772
rect 9306 5692 9312 5704
rect 8036 5664 8248 5692
rect 8496 5664 9312 5692
rect 7616 5596 7788 5624
rect 8205 5627 8263 5633
rect 7616 5584 7622 5596
rect 8205 5593 8217 5627
rect 8251 5624 8263 5627
rect 8496 5624 8524 5664
rect 9306 5652 9312 5664
rect 9364 5692 9370 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9364 5664 9781 5692
rect 9364 5652 9370 5664
rect 9769 5661 9781 5664
rect 9815 5692 9827 5695
rect 9968 5692 9996 5800
rect 14918 5788 14924 5800
rect 14976 5788 14982 5840
rect 11974 5720 11980 5772
rect 12032 5720 12038 5772
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 9815 5664 9996 5692
rect 12084 5688 12112 5723
rect 9815 5661 9827 5664
rect 9769 5655 9827 5661
rect 11992 5660 12112 5688
rect 8251 5596 8524 5624
rect 8573 5627 8631 5633
rect 8251 5593 8263 5596
rect 8205 5587 8263 5593
rect 8573 5593 8585 5627
rect 8619 5624 8631 5627
rect 8938 5624 8944 5636
rect 8619 5596 8944 5624
rect 8619 5593 8631 5596
rect 8573 5587 8631 5593
rect 8938 5584 8944 5596
rect 8996 5624 9002 5636
rect 11882 5624 11888 5636
rect 8996 5596 11888 5624
rect 8996 5584 9002 5596
rect 11882 5584 11888 5596
rect 11940 5584 11946 5636
rect 11992 5624 12020 5660
rect 12158 5652 12164 5704
rect 12216 5652 12222 5704
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 12618 5692 12624 5704
rect 12299 5664 12624 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5692 15531 5695
rect 18138 5692 18144 5704
rect 15519 5664 18144 5692
rect 15519 5661 15531 5664
rect 15473 5655 15531 5661
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 13998 5624 14004 5636
rect 11992 5596 14004 5624
rect 13998 5584 14004 5596
rect 14056 5624 14062 5636
rect 18414 5624 18420 5636
rect 14056 5596 18420 5624
rect 14056 5584 14062 5596
rect 18414 5584 18420 5596
rect 18472 5584 18478 5636
rect 4172 5528 7144 5556
rect 7193 5559 7251 5565
rect 1544 5516 1550 5528
rect 7193 5525 7205 5559
rect 7239 5556 7251 5559
rect 8110 5556 8116 5568
rect 7239 5528 8116 5556
rect 7239 5525 7251 5528
rect 7193 5519 7251 5525
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8294 5516 8300 5568
rect 8352 5516 8358 5568
rect 8389 5559 8447 5565
rect 8389 5525 8401 5559
rect 8435 5556 8447 5559
rect 8754 5556 8760 5568
rect 8435 5528 8760 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 9214 5516 9220 5568
rect 9272 5556 9278 5568
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 9272 5528 11805 5556
rect 9272 5516 9278 5528
rect 11793 5525 11805 5528
rect 11839 5525 11851 5559
rect 11793 5519 11851 5525
rect 16850 5516 16856 5568
rect 16908 5556 16914 5568
rect 18046 5556 18052 5568
rect 16908 5528 18052 5556
rect 16908 5516 16914 5528
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 1104 5466 18860 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 17610 5466
rect 17662 5414 17674 5466
rect 17726 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 18860 5466
rect 1104 5392 18860 5414
rect 1857 5355 1915 5361
rect 1857 5321 1869 5355
rect 1903 5352 1915 5355
rect 10042 5352 10048 5364
rect 1903 5324 10048 5352
rect 1903 5321 1915 5324
rect 1857 5315 1915 5321
rect 10042 5312 10048 5324
rect 10100 5352 10106 5364
rect 10870 5352 10876 5364
rect 10100 5324 10876 5352
rect 10100 5312 10106 5324
rect 10870 5312 10876 5324
rect 10928 5312 10934 5364
rect 11701 5355 11759 5361
rect 11701 5321 11713 5355
rect 11747 5352 11759 5355
rect 14182 5352 14188 5364
rect 11747 5324 14188 5352
rect 11747 5321 11759 5324
rect 11701 5315 11759 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 15010 5312 15016 5364
rect 15068 5352 15074 5364
rect 15841 5355 15899 5361
rect 15841 5352 15853 5355
rect 15068 5324 15853 5352
rect 15068 5312 15074 5324
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 3878 5284 3884 5296
rect 1811 5256 3884 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 3970 5244 3976 5296
rect 4028 5244 4034 5296
rect 5442 5284 5448 5296
rect 5198 5256 5448 5284
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 6362 5244 6368 5296
rect 6420 5284 6426 5296
rect 6822 5284 6828 5296
rect 6420 5256 6828 5284
rect 6420 5244 6426 5256
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 7650 5284 7656 5296
rect 7392 5256 7656 5284
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 3142 5216 3148 5228
rect 2455 5188 3148 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 3697 5219 3755 5225
rect 3697 5216 3709 5219
rect 3660 5188 3709 5216
rect 3660 5176 3666 5188
rect 3697 5185 3709 5188
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 6546 5176 6552 5228
rect 6604 5216 6610 5228
rect 7392 5216 7420 5256
rect 7650 5244 7656 5256
rect 7708 5244 7714 5296
rect 7837 5287 7895 5293
rect 7837 5253 7849 5287
rect 7883 5284 7895 5287
rect 9766 5284 9772 5296
rect 7883 5256 9772 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 9766 5244 9772 5256
rect 9824 5244 9830 5296
rect 11606 5244 11612 5296
rect 11664 5284 11670 5296
rect 12253 5287 12311 5293
rect 12253 5284 12265 5287
rect 11664 5256 12265 5284
rect 11664 5244 11670 5256
rect 12253 5253 12265 5256
rect 12299 5253 12311 5287
rect 12253 5247 12311 5253
rect 6604 5188 7420 5216
rect 7469 5219 7527 5225
rect 6604 5176 6610 5188
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 8110 5216 8116 5228
rect 7607 5188 8116 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 2038 5108 2044 5160
rect 2096 5108 2102 5160
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 2547 5120 3832 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 1394 4972 1400 5024
rect 1452 4972 1458 5024
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 1728 4984 2789 5012
rect 1728 4972 1734 4984
rect 2777 4981 2789 4984
rect 2823 4981 2835 5015
rect 3804 5012 3832 5120
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 4028 5120 5457 5148
rect 4028 5108 4034 5120
rect 5445 5117 5457 5120
rect 5491 5148 5503 5151
rect 6270 5148 6276 5160
rect 5491 5120 6276 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 7484 5148 7512 5179
rect 8110 5176 8116 5188
rect 8168 5216 8174 5228
rect 9582 5216 9588 5228
rect 8168 5188 9588 5216
rect 8168 5176 8174 5188
rect 9582 5176 9588 5188
rect 9640 5216 9646 5228
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 9640 5188 11805 5216
rect 9640 5176 9646 5188
rect 11793 5185 11805 5188
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 11882 5176 11888 5228
rect 11940 5176 11946 5228
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5216 12219 5219
rect 12342 5216 12348 5228
rect 12207 5188 12348 5216
rect 12207 5185 12219 5188
rect 12161 5179 12219 5185
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 15672 5216 15700 5324
rect 15841 5321 15853 5324
rect 15887 5321 15899 5355
rect 15841 5315 15899 5321
rect 15749 5287 15807 5293
rect 15749 5253 15761 5287
rect 15795 5284 15807 5287
rect 18322 5284 18328 5296
rect 15795 5256 18328 5284
rect 15795 5253 15807 5256
rect 15749 5247 15807 5253
rect 18322 5244 18328 5256
rect 18380 5244 18386 5296
rect 16025 5219 16083 5225
rect 16025 5216 16037 5219
rect 15672 5188 16037 5216
rect 16025 5185 16037 5188
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 8478 5148 8484 5160
rect 6420 5120 8484 5148
rect 6420 5108 6426 5120
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 9950 5148 9956 5160
rect 9824 5120 9956 5148
rect 9824 5108 9830 5120
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 12066 5148 12072 5160
rect 10192 5120 12072 5148
rect 10192 5108 10198 5120
rect 12066 5108 12072 5120
rect 12124 5108 12130 5160
rect 7282 5040 7288 5092
rect 7340 5040 7346 5092
rect 10962 5040 10968 5092
rect 11020 5080 11026 5092
rect 11517 5083 11575 5089
rect 11517 5080 11529 5083
rect 11020 5052 11529 5080
rect 11020 5040 11026 5052
rect 11517 5049 11529 5052
rect 11563 5049 11575 5083
rect 11517 5043 11575 5049
rect 15194 5040 15200 5092
rect 15252 5080 15258 5092
rect 16209 5083 16267 5089
rect 16209 5080 16221 5083
rect 15252 5052 16221 5080
rect 15252 5040 15258 5052
rect 16209 5049 16221 5052
rect 16255 5049 16267 5083
rect 16209 5043 16267 5049
rect 5442 5012 5448 5024
rect 3804 4984 5448 5012
rect 2777 4975 2835 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 10226 4972 10232 5024
rect 10284 5012 10290 5024
rect 11698 5012 11704 5024
rect 10284 4984 11704 5012
rect 10284 4972 10290 4984
rect 11698 4972 11704 4984
rect 11756 5012 11762 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 11756 4984 12081 5012
rect 11756 4972 11762 4984
rect 12069 4981 12081 4984
rect 12115 4981 12127 5015
rect 12069 4975 12127 4981
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 17862 5012 17868 5024
rect 17460 4984 17868 5012
rect 17460 4972 17466 4984
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 1104 4922 18860 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 16950 4922
rect 17002 4870 17014 4922
rect 17066 4870 17078 4922
rect 17130 4870 17142 4922
rect 17194 4870 17206 4922
rect 17258 4870 18860 4922
rect 1104 4848 18860 4870
rect 1412 4780 3096 4808
rect 1412 4681 1440 4780
rect 3068 4740 3096 4780
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 5258 4768 5264 4820
rect 5316 4768 5322 4820
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4808 7435 4811
rect 7650 4808 7656 4820
rect 7423 4780 7656 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 9490 4768 9496 4820
rect 9548 4808 9554 4820
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 9548 4780 9597 4808
rect 9548 4768 9554 4780
rect 9585 4777 9597 4780
rect 9631 4777 9643 4811
rect 16850 4808 16856 4820
rect 9585 4771 9643 4777
rect 9692 4780 16856 4808
rect 3602 4740 3608 4752
rect 3068 4712 3608 4740
rect 3602 4700 3608 4712
rect 3660 4700 3666 4752
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 9692 4740 9720 4780
rect 16850 4768 16856 4780
rect 16908 4808 16914 4820
rect 16945 4811 17003 4817
rect 16945 4808 16957 4811
rect 16908 4780 16957 4808
rect 16908 4768 16914 4780
rect 16945 4777 16957 4780
rect 16991 4808 17003 4811
rect 17402 4808 17408 4820
rect 16991 4780 17408 4808
rect 16991 4777 17003 4780
rect 16945 4771 17003 4777
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 10410 4740 10416 4752
rect 7340 4712 9720 4740
rect 9784 4712 10416 4740
rect 7340 4700 7346 4712
rect 4988 4684 5040 4690
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4641 1455 4675
rect 1397 4635 1455 4641
rect 1670 4632 1676 4684
rect 1728 4632 1734 4684
rect 5902 4672 5908 4684
rect 5040 4644 5908 4672
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 6012 4644 7420 4672
rect 4988 4626 5040 4632
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 6012 4613 6040 4644
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 6696 4576 6745 4604
rect 6696 4564 6702 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6972 4576 7021 4604
rect 6972 4564 6978 4576
rect 7009 4573 7021 4576
rect 7055 4604 7067 4607
rect 7190 4604 7196 4616
rect 7055 4576 7196 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 7392 4604 7420 4644
rect 7466 4632 7472 4684
rect 7524 4672 7530 4684
rect 9674 4672 9680 4684
rect 7524 4644 9680 4672
rect 7524 4632 7530 4644
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9784 4672 9812 4712
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 9784 4644 9904 4672
rect 7392 4576 9720 4604
rect 3050 4536 3056 4548
rect 2898 4508 3056 4536
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 3418 4496 3424 4548
rect 3476 4536 3482 4548
rect 3973 4539 4031 4545
rect 3973 4536 3985 4539
rect 3476 4508 3985 4536
rect 3476 4496 3482 4508
rect 3973 4505 3985 4508
rect 4019 4505 4031 4539
rect 3973 4499 4031 4505
rect 4341 4539 4399 4545
rect 4341 4505 4353 4539
rect 4387 4536 4399 4539
rect 4522 4536 4528 4548
rect 4387 4508 4528 4536
rect 4387 4505 4399 4508
rect 4341 4499 4399 4505
rect 2038 4428 2044 4480
rect 2096 4468 2102 4480
rect 4356 4468 4384 4499
rect 4522 4496 4528 4508
rect 4580 4496 4586 4548
rect 4709 4539 4767 4545
rect 4709 4505 4721 4539
rect 4755 4536 4767 4539
rect 5350 4536 5356 4548
rect 4755 4508 5356 4536
rect 4755 4505 4767 4508
rect 4709 4499 4767 4505
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 6822 4496 6828 4548
rect 6880 4536 6886 4548
rect 9692 4536 9720 4576
rect 9766 4564 9772 4616
rect 9824 4564 9830 4616
rect 9876 4613 9904 4644
rect 10042 4632 10048 4684
rect 10100 4632 10106 4684
rect 11882 4632 11888 4684
rect 11940 4632 11946 4684
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 12032 4644 13768 4672
rect 12032 4632 12038 4644
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10008 4576 10053 4604
rect 10008 4564 10014 4576
rect 11422 4564 11428 4616
rect 11480 4604 11486 4616
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11480 4576 11621 4604
rect 11480 4564 11486 4576
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 13740 4604 13768 4644
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 13872 4644 15485 4672
rect 13872 4632 13878 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 15473 4635 15531 4641
rect 15194 4604 15200 4616
rect 13740 4576 15200 4604
rect 11609 4567 11667 4573
rect 10318 4536 10324 4548
rect 6880 4508 7604 4536
rect 9692 4508 10324 4536
rect 6880 4496 6886 4508
rect 2096 4440 4384 4468
rect 2096 4428 2102 4440
rect 4430 4428 4436 4480
rect 4488 4468 4494 4480
rect 5077 4471 5135 4477
rect 5077 4468 5089 4471
rect 4488 4440 5089 4468
rect 4488 4428 4494 4440
rect 5077 4437 5089 4440
rect 5123 4437 5135 4471
rect 5077 4431 5135 4437
rect 7374 4428 7380 4480
rect 7432 4428 7438 4480
rect 7576 4477 7604 4508
rect 10318 4496 10324 4508
rect 10376 4496 10382 4548
rect 11624 4536 11652 4567
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 11790 4536 11796 4548
rect 11624 4508 11796 4536
rect 11790 4496 11796 4508
rect 11848 4536 11854 4548
rect 11974 4536 11980 4548
rect 11848 4508 11980 4536
rect 11848 4496 11854 4508
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 12526 4496 12532 4548
rect 12584 4496 12590 4548
rect 15746 4496 15752 4548
rect 15804 4536 15810 4548
rect 15804 4508 15962 4536
rect 15804 4496 15810 4508
rect 7561 4471 7619 4477
rect 7561 4437 7573 4471
rect 7607 4437 7619 4471
rect 7561 4431 7619 4437
rect 8018 4428 8024 4480
rect 8076 4468 8082 4480
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 8076 4440 13369 4468
rect 8076 4428 8082 4440
rect 13357 4437 13369 4440
rect 13403 4437 13415 4471
rect 13357 4431 13415 4437
rect 1104 4378 18860 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 17610 4378
rect 17662 4326 17674 4378
rect 17726 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 18860 4378
rect 1104 4304 18860 4326
rect 2343 4267 2401 4273
rect 2343 4233 2355 4267
rect 2389 4264 2401 4267
rect 3326 4264 3332 4276
rect 2389 4236 3332 4264
rect 2389 4233 2401 4236
rect 2343 4227 2401 4233
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 5813 4267 5871 4273
rect 5813 4233 5825 4267
rect 5859 4233 5871 4267
rect 5813 4227 5871 4233
rect 2130 4156 2136 4208
rect 2188 4156 2194 4208
rect 4798 4156 4804 4208
rect 4856 4156 4862 4208
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4128 1547 4131
rect 1578 4128 1584 4140
rect 1535 4100 1584 4128
rect 1535 4097 1547 4100
rect 1489 4091 1547 4097
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 1670 4088 1676 4140
rect 1728 4088 1734 4140
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4128 2007 4131
rect 2222 4128 2228 4140
rect 1995 4100 2228 4128
rect 1995 4097 2007 4100
rect 1949 4091 2007 4097
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 3602 4088 3608 4140
rect 3660 4128 3666 4140
rect 4065 4131 4123 4137
rect 4065 4128 4077 4131
rect 3660 4100 4077 4128
rect 3660 4088 3666 4100
rect 4065 4097 4077 4100
rect 4111 4097 4123 4131
rect 5828 4128 5856 4227
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 14182 4264 14188 4276
rect 8536 4236 14188 4264
rect 8536 4224 8542 4236
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 17494 4224 17500 4276
rect 17552 4264 17558 4276
rect 18233 4267 18291 4273
rect 18233 4264 18245 4267
rect 17552 4236 18245 4264
rect 17552 4224 17558 4236
rect 18233 4233 18245 4236
rect 18279 4233 18291 4267
rect 18233 4227 18291 4233
rect 18414 4224 18420 4276
rect 18472 4224 18478 4276
rect 8386 4196 8392 4208
rect 7024 4168 7512 4196
rect 7024 4128 7052 4168
rect 5828 4100 7052 4128
rect 7116 4100 7420 4128
rect 4065 4091 4123 4097
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4060 1823 4063
rect 3878 4060 3884 4072
rect 1811 4032 3884 4060
rect 1811 4029 1823 4032
rect 1765 4023 1823 4029
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4060 4399 4063
rect 7116 4060 7144 4100
rect 4387 4032 7144 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 1857 3995 1915 4001
rect 1857 3961 1869 3995
rect 1903 3992 1915 3995
rect 2038 3992 2044 4004
rect 1903 3964 2044 3992
rect 1903 3961 1915 3964
rect 1857 3955 1915 3961
rect 2038 3952 2044 3964
rect 2096 3952 2102 4004
rect 2498 3952 2504 4004
rect 2556 3952 2562 4004
rect 7392 3992 7420 4100
rect 7484 4060 7512 4168
rect 8128 4168 8392 4196
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4128 7619 4131
rect 8128 4128 8156 4168
rect 8386 4156 8392 4168
rect 8444 4156 8450 4208
rect 13262 4196 13268 4208
rect 13018 4168 13268 4196
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 14550 4156 14556 4208
rect 14608 4196 14614 4208
rect 18046 4196 18052 4208
rect 14608 4168 18052 4196
rect 14608 4156 14614 4168
rect 18046 4156 18052 4168
rect 18104 4156 18110 4208
rect 7607 4100 8156 4128
rect 8205 4131 8263 4137
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 8205 4097 8217 4131
rect 8251 4128 8263 4131
rect 9950 4128 9956 4140
rect 8251 4100 9956 4128
rect 8251 4097 8263 4100
rect 8205 4091 8263 4097
rect 8220 4060 8248 4091
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 13004 4100 16681 4128
rect 7484 4032 8248 4060
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8478 4060 8484 4072
rect 8343 4032 8484 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 11422 4060 11428 4072
rect 8996 4032 11428 4060
rect 8996 4020 9002 4032
rect 11422 4020 11428 4032
rect 11480 4060 11486 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11480 4032 11529 4060
rect 11480 4020 11486 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11517 4023 11575 4029
rect 11790 4020 11796 4072
rect 11848 4020 11854 4072
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 13004 4060 13032 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 11940 4032 13032 4060
rect 11940 4020 11946 4032
rect 14182 4020 14188 4072
rect 14240 4060 14246 4072
rect 14240 4032 17540 4060
rect 14240 4020 14246 4032
rect 8573 3995 8631 4001
rect 8573 3992 8585 3995
rect 7392 3964 8585 3992
rect 8573 3961 8585 3964
rect 8619 3961 8631 3995
rect 8573 3955 8631 3961
rect 15654 3952 15660 4004
rect 15712 3992 15718 4004
rect 16945 3995 17003 4001
rect 16945 3992 16957 3995
rect 15712 3964 16957 3992
rect 15712 3952 15718 3964
rect 16945 3961 16957 3964
rect 16991 3992 17003 3995
rect 17405 3995 17463 4001
rect 17405 3992 17417 3995
rect 16991 3964 17417 3992
rect 16991 3961 17003 3964
rect 16945 3955 17003 3961
rect 17405 3961 17417 3964
rect 17451 3961 17463 3995
rect 17512 3992 17540 4032
rect 17586 4020 17592 4072
rect 17644 4060 17650 4072
rect 18690 4060 18696 4072
rect 17644 4032 18696 4060
rect 17644 4020 17650 4032
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 18138 3992 18144 4004
rect 17512 3964 18144 3992
rect 17405 3955 17463 3961
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 3050 3924 3056 3936
rect 2363 3896 3056 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 5074 3924 5080 3936
rect 4396 3896 5080 3924
rect 4396 3884 4402 3896
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 7377 3927 7435 3933
rect 7377 3893 7389 3927
rect 7423 3924 7435 3927
rect 9582 3924 9588 3936
rect 7423 3896 9588 3924
rect 7423 3893 7435 3896
rect 7377 3887 7435 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 13265 3927 13323 3933
rect 13265 3924 13277 3927
rect 9732 3896 13277 3924
rect 9732 3884 9738 3896
rect 13265 3893 13277 3896
rect 13311 3893 13323 3927
rect 13265 3887 13323 3893
rect 15286 3884 15292 3936
rect 15344 3924 15350 3936
rect 17129 3927 17187 3933
rect 17129 3924 17141 3927
rect 15344 3896 17141 3924
rect 15344 3884 15350 3896
rect 17129 3893 17141 3896
rect 17175 3893 17187 3927
rect 17129 3887 17187 3893
rect 18233 3927 18291 3933
rect 18233 3893 18245 3927
rect 18279 3924 18291 3927
rect 18598 3924 18604 3936
rect 18279 3896 18604 3924
rect 18279 3893 18291 3896
rect 18233 3887 18291 3893
rect 18598 3884 18604 3896
rect 18656 3884 18662 3936
rect 1104 3834 18860 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 16950 3834
rect 17002 3782 17014 3834
rect 17066 3782 17078 3834
rect 17130 3782 17142 3834
rect 17194 3782 17206 3834
rect 17258 3782 18860 3834
rect 1104 3760 18860 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 1854 3720 1860 3732
rect 1627 3692 1860 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 4617 3723 4675 3729
rect 4617 3689 4629 3723
rect 4663 3720 4675 3723
rect 5534 3720 5540 3732
rect 4663 3692 5540 3720
rect 4663 3689 4675 3692
rect 4617 3683 4675 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 9674 3720 9680 3732
rect 6512 3692 9680 3720
rect 6512 3680 6518 3692
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 14810 3723 14868 3729
rect 14810 3720 14822 3723
rect 11112 3692 14822 3720
rect 11112 3680 11118 3692
rect 14810 3689 14822 3692
rect 14856 3720 14868 3723
rect 14856 3692 16804 3720
rect 14856 3689 14868 3692
rect 14810 3683 14868 3689
rect 1489 3655 1547 3661
rect 1489 3621 1501 3655
rect 1535 3652 1547 3655
rect 3694 3652 3700 3664
rect 1535 3624 3700 3652
rect 1535 3621 1547 3624
rect 1489 3615 1547 3621
rect 3694 3612 3700 3624
rect 3752 3612 3758 3664
rect 3881 3655 3939 3661
rect 3881 3621 3893 3655
rect 3927 3652 3939 3655
rect 4246 3652 4252 3664
rect 3927 3624 4252 3652
rect 3927 3621 3939 3624
rect 3881 3615 3939 3621
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 4890 3652 4896 3664
rect 4448 3624 4896 3652
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 2314 3584 2320 3596
rect 1719 3556 2320 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 4338 3584 4344 3596
rect 2746 3556 4344 3584
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3516 1823 3519
rect 2746 3516 2774 3556
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 4448 3593 4476 3624
rect 4890 3612 4896 3624
rect 4948 3652 4954 3664
rect 4948 3624 5764 3652
rect 4948 3612 4954 3624
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3553 4491 3587
rect 4433 3547 4491 3553
rect 5442 3544 5448 3596
rect 5500 3544 5506 3596
rect 5736 3584 5764 3624
rect 5810 3612 5816 3664
rect 5868 3612 5874 3664
rect 11146 3612 11152 3664
rect 11204 3612 11210 3664
rect 11330 3612 11336 3664
rect 11388 3652 11394 3664
rect 11388 3624 11836 3652
rect 11388 3612 11394 3624
rect 7374 3584 7380 3596
rect 5736 3556 7380 3584
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 9306 3544 9312 3596
rect 9364 3584 9370 3596
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 9364 3556 10977 3584
rect 9364 3544 9370 3556
rect 10965 3553 10977 3556
rect 11011 3584 11023 3587
rect 11698 3584 11704 3596
rect 11011 3556 11704 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 11808 3593 11836 3624
rect 14550 3612 14556 3664
rect 14608 3652 14614 3664
rect 14921 3655 14979 3661
rect 14921 3652 14933 3655
rect 14608 3624 14933 3652
rect 14608 3612 14614 3624
rect 14921 3621 14933 3624
rect 14967 3621 14979 3655
rect 16776 3652 16804 3692
rect 17494 3680 17500 3732
rect 17552 3680 17558 3732
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 18233 3723 18291 3729
rect 18233 3720 18245 3723
rect 18196 3692 18245 3720
rect 18196 3680 18202 3692
rect 18233 3689 18245 3692
rect 18279 3689 18291 3723
rect 18233 3683 18291 3689
rect 18598 3652 18604 3664
rect 14921 3615 14979 3621
rect 15028 3624 15608 3652
rect 16776 3624 18604 3652
rect 11793 3587 11851 3593
rect 11793 3553 11805 3587
rect 11839 3553 11851 3587
rect 11793 3547 11851 3553
rect 12158 3544 12164 3596
rect 12216 3584 12222 3596
rect 15028 3593 15056 3624
rect 15013 3587 15071 3593
rect 15013 3584 15025 3587
rect 12216 3556 15025 3584
rect 12216 3544 12222 3556
rect 15013 3553 15025 3556
rect 15059 3553 15071 3587
rect 15013 3547 15071 3553
rect 15102 3544 15108 3596
rect 15160 3544 15166 3596
rect 15194 3544 15200 3596
rect 15252 3584 15258 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 15252 3556 15485 3584
rect 15252 3544 15258 3556
rect 15473 3553 15485 3556
rect 15519 3553 15531 3587
rect 15580 3584 15608 3624
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 18506 3584 18512 3596
rect 15580 3556 18512 3584
rect 15473 3547 15531 3553
rect 18506 3544 18512 3556
rect 18564 3544 18570 3596
rect 7282 3516 7288 3528
rect 1811 3488 2774 3516
rect 4264 3488 7288 3516
rect 1811 3485 1823 3488
rect 1765 3479 1823 3485
rect 1412 3448 1440 3479
rect 1412 3420 1900 3448
rect 1872 3392 1900 3420
rect 3878 3408 3884 3460
rect 3936 3448 3942 3460
rect 4264 3448 4292 3488
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 8938 3476 8944 3528
rect 8996 3476 9002 3528
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 3936 3420 4292 3448
rect 4341 3451 4399 3457
rect 3936 3408 3942 3420
rect 4341 3417 4353 3451
rect 4387 3448 4399 3451
rect 4522 3448 4528 3460
rect 4387 3420 4528 3448
rect 4387 3417 4399 3420
rect 4341 3411 4399 3417
rect 4522 3408 4528 3420
rect 4580 3448 4586 3460
rect 8846 3448 8852 3460
rect 4580 3420 8852 3448
rect 4580 3408 4586 3420
rect 8846 3408 8852 3420
rect 8904 3448 8910 3460
rect 9122 3448 9128 3460
rect 8904 3420 9128 3448
rect 8904 3408 8910 3420
rect 9122 3408 9128 3420
rect 9180 3408 9186 3460
rect 9214 3408 9220 3460
rect 9272 3408 9278 3460
rect 10870 3448 10876 3460
rect 10442 3420 10876 3448
rect 10870 3408 10876 3420
rect 10928 3408 10934 3460
rect 1854 3340 1860 3392
rect 1912 3340 1918 3392
rect 5905 3383 5963 3389
rect 5905 3349 5917 3383
rect 5951 3380 5963 3383
rect 9490 3380 9496 3392
rect 5951 3352 9496 3380
rect 5951 3349 5963 3352
rect 5905 3343 5963 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 11072 3380 11100 3479
rect 11882 3476 11888 3528
rect 11940 3476 11946 3528
rect 12250 3476 12256 3528
rect 12308 3476 12314 3528
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 13170 3516 13176 3528
rect 12575 3488 13176 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 13596 3488 14657 3516
rect 13596 3476 13602 3488
rect 14645 3485 14657 3488
rect 14691 3485 14703 3519
rect 14645 3479 14703 3485
rect 17405 3519 17463 3525
rect 17405 3485 17417 3519
rect 17451 3516 17463 3519
rect 17862 3516 17868 3528
rect 17451 3488 17868 3516
rect 17451 3485 17463 3488
rect 17405 3479 17463 3485
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 12066 3408 12072 3460
rect 12124 3448 12130 3460
rect 15654 3448 15660 3460
rect 12124 3420 15660 3448
rect 12124 3408 12130 3420
rect 15654 3408 15660 3420
rect 15712 3408 15718 3460
rect 15746 3408 15752 3460
rect 15804 3408 15810 3460
rect 17310 3448 17316 3460
rect 16974 3420 17316 3448
rect 17310 3408 17316 3420
rect 17368 3408 17374 3460
rect 18138 3408 18144 3460
rect 18196 3408 18202 3460
rect 9640 3352 11100 3380
rect 9640 3340 9646 3352
rect 14642 3340 14648 3392
rect 14700 3380 14706 3392
rect 17221 3383 17279 3389
rect 17221 3380 17233 3383
rect 14700 3352 17233 3380
rect 14700 3340 14706 3352
rect 17221 3349 17233 3352
rect 17267 3349 17279 3383
rect 17221 3343 17279 3349
rect 1104 3290 18860 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 17610 3290
rect 17662 3238 17674 3290
rect 17726 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 18860 3290
rect 1104 3216 18860 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 6086 3176 6092 3188
rect 1912 3148 6092 3176
rect 1912 3136 1918 3148
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6196 3148 6500 3176
rect 1489 3111 1547 3117
rect 1489 3077 1501 3111
rect 1535 3108 1547 3111
rect 3050 3108 3056 3120
rect 1535 3080 3056 3108
rect 1535 3077 1547 3080
rect 1489 3071 1547 3077
rect 3050 3068 3056 3080
rect 3108 3108 3114 3120
rect 4062 3108 4068 3120
rect 3108 3080 4068 3108
rect 3108 3068 3114 3080
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 6196 3108 6224 3148
rect 5500 3080 6224 3108
rect 5500 3068 5506 3080
rect 6362 3068 6368 3120
rect 6420 3068 6426 3120
rect 6472 3108 6500 3148
rect 6546 3136 6552 3188
rect 6604 3185 6610 3188
rect 6604 3179 6623 3185
rect 6611 3145 6623 3179
rect 6604 3139 6623 3145
rect 6733 3179 6791 3185
rect 6733 3145 6745 3179
rect 6779 3145 6791 3179
rect 9582 3176 9588 3188
rect 6733 3139 6791 3145
rect 9048 3148 9588 3176
rect 6604 3136 6610 3139
rect 6748 3108 6776 3139
rect 6472 3080 6776 3108
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 4246 3040 4252 3052
rect 1728 3012 4252 3040
rect 1728 3000 1734 3012
rect 4246 3000 4252 3012
rect 4304 3040 4310 3052
rect 9048 3040 9076 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9677 3179 9735 3185
rect 9677 3145 9689 3179
rect 9723 3176 9735 3179
rect 9858 3176 9864 3188
rect 9723 3148 9864 3176
rect 9723 3145 9735 3148
rect 9677 3139 9735 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10505 3179 10563 3185
rect 10505 3145 10517 3179
rect 10551 3176 10563 3179
rect 12250 3176 12256 3188
rect 10551 3148 12256 3176
rect 10551 3145 10563 3148
rect 10505 3139 10563 3145
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 13173 3179 13231 3185
rect 13173 3145 13185 3179
rect 13219 3176 13231 3179
rect 13354 3176 13360 3188
rect 13219 3148 13360 3176
rect 13219 3145 13231 3148
rect 13173 3139 13231 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 16317 3179 16375 3185
rect 16317 3176 16329 3179
rect 15436 3148 16329 3176
rect 15436 3136 15442 3148
rect 16317 3145 16329 3148
rect 16363 3145 16375 3179
rect 16317 3139 16375 3145
rect 16482 3136 16488 3188
rect 16540 3136 16546 3188
rect 9122 3068 9128 3120
rect 9180 3108 9186 3120
rect 11054 3108 11060 3120
rect 9180 3080 11060 3108
rect 9180 3068 9186 3080
rect 4304 3012 9076 3040
rect 4304 3000 4310 3012
rect 9490 3000 9496 3052
rect 9548 3000 9554 3052
rect 10704 3049 10732 3080
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 14550 3108 14556 3120
rect 11204 3080 14556 3108
rect 11204 3068 11210 3080
rect 14550 3068 14556 3080
rect 14608 3068 14614 3120
rect 14918 3068 14924 3120
rect 14976 3108 14982 3120
rect 16117 3111 16175 3117
rect 16117 3108 16129 3111
rect 14976 3080 16129 3108
rect 14976 3068 14982 3080
rect 16117 3077 16129 3080
rect 16163 3108 16175 3111
rect 17586 3108 17592 3120
rect 16163 3080 17592 3108
rect 16163 3077 16175 3080
rect 16117 3071 16175 3077
rect 17586 3068 17592 3080
rect 17644 3068 17650 3120
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3040 11023 3043
rect 11514 3040 11520 3052
rect 11011 3012 11520 3040
rect 11011 3009 11023 3012
rect 10965 3003 11023 3009
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11756 3012 12434 3040
rect 11756 3000 11762 3012
rect 4062 2932 4068 2984
rect 4120 2972 4126 2984
rect 11330 2972 11336 2984
rect 4120 2944 11336 2972
rect 4120 2932 4126 2944
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 11606 2932 11612 2984
rect 11664 2932 11670 2984
rect 12406 2972 12434 3012
rect 13078 3000 13084 3052
rect 13136 3000 13142 3052
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14240 3012 14841 3040
rect 14240 3000 14246 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 15286 3000 15292 3052
rect 15344 3000 15350 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 17129 3043 17187 3049
rect 17129 3040 17141 3043
rect 16816 3012 17141 3040
rect 16816 3000 16822 3012
rect 17129 3009 17141 3012
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 17402 3000 17408 3052
rect 17460 3000 17466 3052
rect 16206 2972 16212 2984
rect 12406 2944 16212 2972
rect 16206 2932 16212 2944
rect 16264 2932 16270 2984
rect 16298 2932 16304 2984
rect 16356 2972 16362 2984
rect 16945 2975 17003 2981
rect 16945 2972 16957 2975
rect 16356 2944 16957 2972
rect 16356 2932 16362 2944
rect 16945 2941 16957 2944
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2972 17371 2975
rect 18782 2972 18788 2984
rect 17359 2944 18788 2972
rect 17359 2941 17371 2944
rect 17313 2935 17371 2941
rect 8110 2904 8116 2916
rect 6555 2876 8116 2904
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 6555 2845 6583 2876
rect 8110 2864 8116 2876
rect 8168 2864 8174 2916
rect 9214 2864 9220 2916
rect 9272 2904 9278 2916
rect 12069 2907 12127 2913
rect 12069 2904 12081 2907
rect 9272 2876 12081 2904
rect 9272 2864 9278 2876
rect 12069 2873 12081 2876
rect 12115 2873 12127 2907
rect 12069 2867 12127 2873
rect 12986 2864 12992 2916
rect 13044 2904 13050 2916
rect 13044 2876 14044 2904
rect 13044 2864 13050 2876
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 992 2808 1593 2836
rect 992 2796 998 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 6549 2839 6607 2845
rect 6549 2805 6561 2839
rect 6595 2805 6607 2839
rect 6549 2799 6607 2805
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 10873 2839 10931 2845
rect 10873 2836 10885 2839
rect 7340 2808 10885 2836
rect 7340 2796 7346 2808
rect 10873 2805 10885 2808
rect 10919 2836 10931 2839
rect 11146 2836 11152 2848
rect 10919 2808 11152 2836
rect 10919 2805 10931 2808
rect 10873 2799 10931 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11330 2796 11336 2848
rect 11388 2836 11394 2848
rect 13906 2836 13912 2848
rect 11388 2808 13912 2836
rect 11388 2796 11394 2808
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 14016 2836 14044 2876
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 15473 2907 15531 2913
rect 15473 2904 15485 2907
rect 14884 2876 15485 2904
rect 14884 2864 14890 2876
rect 15473 2873 15485 2876
rect 15519 2873 15531 2907
rect 17236 2904 17264 2935
rect 17494 2904 17500 2916
rect 15473 2867 15531 2873
rect 16040 2876 16436 2904
rect 17236 2876 17500 2904
rect 15105 2839 15163 2845
rect 15105 2836 15117 2839
rect 14016 2808 15117 2836
rect 15105 2805 15117 2808
rect 15151 2836 15163 2839
rect 16040 2836 16068 2876
rect 15151 2808 16068 2836
rect 15151 2805 15163 2808
rect 15105 2799 15163 2805
rect 16298 2796 16304 2848
rect 16356 2796 16362 2848
rect 16408 2836 16436 2876
rect 17494 2864 17500 2876
rect 17552 2864 17558 2916
rect 17604 2836 17632 2944
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 16408 2808 17632 2836
rect 1104 2746 18860 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 16950 2746
rect 17002 2694 17014 2746
rect 17066 2694 17078 2746
rect 17130 2694 17142 2746
rect 17194 2694 17206 2746
rect 17258 2694 18860 2746
rect 1104 2672 18860 2694
rect 5902 2592 5908 2644
rect 5960 2632 5966 2644
rect 6089 2635 6147 2641
rect 6089 2632 6101 2635
rect 5960 2604 6101 2632
rect 5960 2592 5966 2604
rect 6089 2601 6101 2604
rect 6135 2601 6147 2635
rect 10962 2632 10968 2644
rect 6089 2595 6147 2601
rect 6886 2604 10968 2632
rect 6178 2496 6184 2508
rect 1504 2468 6184 2496
rect 1504 2437 1532 2468
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 1489 2431 1547 2437
rect 1489 2397 1501 2431
rect 1535 2397 1547 2431
rect 1489 2391 1547 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5868 2400 5917 2428
rect 5868 2388 5874 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 2777 2363 2835 2369
rect 2777 2329 2789 2363
rect 2823 2360 2835 2363
rect 6886 2360 6914 2604
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 13630 2632 13636 2644
rect 11931 2604 13636 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 18322 2592 18328 2644
rect 18380 2592 18386 2644
rect 9122 2524 9128 2576
rect 9180 2524 9186 2576
rect 11790 2524 11796 2576
rect 11848 2564 11854 2576
rect 16298 2564 16304 2576
rect 11848 2536 16304 2564
rect 11848 2524 11854 2536
rect 16298 2524 16304 2536
rect 16356 2524 16362 2576
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 9309 2499 9367 2505
rect 9309 2496 9321 2499
rect 8996 2468 9321 2496
rect 8996 2456 9002 2468
rect 9309 2465 9321 2468
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 10008 2468 14412 2496
rect 10008 2456 10014 2468
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8662 2428 8668 2440
rect 8435 2400 8668 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9033 2431 9091 2437
rect 9033 2397 9045 2431
rect 9079 2428 9091 2431
rect 9079 2400 9260 2428
rect 9079 2397 9091 2400
rect 9033 2391 9091 2397
rect 2823 2332 6914 2360
rect 2823 2329 2835 2332
rect 2777 2323 2835 2329
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 72 2264 1593 2292
rect 72 2252 78 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 2498 2252 2504 2304
rect 2556 2292 2562 2304
rect 2869 2295 2927 2301
rect 2869 2292 2881 2295
rect 2556 2264 2881 2292
rect 2556 2252 2562 2264
rect 2869 2261 2881 2264
rect 2915 2261 2927 2295
rect 2869 2255 2927 2261
rect 8478 2252 8484 2304
rect 8536 2252 8542 2304
rect 9232 2292 9260 2400
rect 11330 2388 11336 2440
rect 11388 2388 11394 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 14384 2437 14412 2468
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 17586 2388 17592 2440
rect 17644 2388 17650 2440
rect 17954 2388 17960 2440
rect 18012 2428 18018 2440
rect 18509 2431 18567 2437
rect 18509 2428 18521 2431
rect 18012 2400 18521 2428
rect 18012 2388 18018 2400
rect 18509 2397 18521 2400
rect 18555 2397 18567 2431
rect 18509 2391 18567 2397
rect 9490 2320 9496 2372
rect 9548 2360 9554 2372
rect 9585 2363 9643 2369
rect 9585 2360 9597 2363
rect 9548 2332 9597 2360
rect 9548 2320 9554 2332
rect 9585 2329 9597 2332
rect 9631 2329 9643 2363
rect 11238 2360 11244 2372
rect 10810 2332 11244 2360
rect 9585 2323 9643 2329
rect 11238 2320 11244 2332
rect 11296 2320 11302 2372
rect 12342 2292 12348 2304
rect 9232 2264 12348 2292
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14461 2295 14519 2301
rect 14461 2292 14473 2295
rect 14240 2264 14473 2292
rect 14240 2252 14246 2264
rect 14461 2261 14473 2264
rect 14507 2261 14519 2295
rect 14461 2255 14519 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 1104 2202 18860 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 17610 2202
rect 17662 2150 17674 2202
rect 17726 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 7610 17382 7662 17434
rect 7674 17382 7726 17434
rect 7738 17382 7790 17434
rect 7802 17382 7854 17434
rect 7866 17382 7918 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 17610 17382 17662 17434
rect 17674 17382 17726 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 664 17212 716 17264
rect 1492 17187 1544 17196
rect 1492 17153 1501 17187
rect 1501 17153 1535 17187
rect 1535 17153 1544 17187
rect 1492 17144 1544 17153
rect 3056 17212 3108 17264
rect 6460 17280 6512 17332
rect 10876 17280 10928 17332
rect 15476 17280 15528 17332
rect 17960 17280 18012 17332
rect 4068 17187 4120 17196
rect 4068 17153 4077 17187
rect 4077 17153 4111 17187
rect 4111 17153 4120 17187
rect 4068 17144 4120 17153
rect 4528 17187 4580 17196
rect 4528 17153 4537 17187
rect 4537 17153 4571 17187
rect 4571 17153 4580 17187
rect 4528 17144 4580 17153
rect 2964 17008 3016 17060
rect 6276 17144 6328 17196
rect 6644 17187 6696 17196
rect 6644 17153 6653 17187
rect 6653 17153 6687 17187
rect 6687 17153 6696 17187
rect 6644 17144 6696 17153
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 6460 17008 6512 17060
rect 4344 16940 4396 16992
rect 4528 16940 4580 16992
rect 9680 17144 9732 17196
rect 12256 17212 12308 17264
rect 14004 17144 14056 17196
rect 15936 17144 15988 17196
rect 16672 17144 16724 17196
rect 8300 17076 8352 17128
rect 14924 17076 14976 17128
rect 15200 17008 15252 17060
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 10416 16940 10468 16992
rect 12808 16940 12860 16992
rect 13544 16940 13596 16992
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 6950 16838 7002 16890
rect 7014 16838 7066 16890
rect 7078 16838 7130 16890
rect 7142 16838 7194 16890
rect 7206 16838 7258 16890
rect 11950 16838 12002 16890
rect 12014 16838 12066 16890
rect 12078 16838 12130 16890
rect 12142 16838 12194 16890
rect 12206 16838 12258 16890
rect 16950 16838 17002 16890
rect 17014 16838 17066 16890
rect 17078 16838 17130 16890
rect 17142 16838 17194 16890
rect 17206 16838 17258 16890
rect 9220 16736 9272 16788
rect 9312 16736 9364 16788
rect 16304 16736 16356 16788
rect 18052 16736 18104 16788
rect 4344 16668 4396 16720
rect 6920 16668 6972 16720
rect 17960 16668 18012 16720
rect 8300 16600 8352 16652
rect 11796 16600 11848 16652
rect 3792 16464 3844 16516
rect 9864 16532 9916 16584
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 11060 16464 11112 16516
rect 12992 16464 13044 16516
rect 17316 16532 17368 16584
rect 16856 16464 16908 16516
rect 10232 16396 10284 16448
rect 13636 16396 13688 16448
rect 16488 16396 16540 16448
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 7610 16294 7662 16346
rect 7674 16294 7726 16346
rect 7738 16294 7790 16346
rect 7802 16294 7854 16346
rect 7866 16294 7918 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 17610 16294 17662 16346
rect 17674 16294 17726 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 6920 16124 6972 16176
rect 3056 16056 3108 16108
rect 3332 16099 3384 16108
rect 3332 16065 3341 16099
rect 3341 16065 3375 16099
rect 3375 16065 3384 16099
rect 3332 16056 3384 16065
rect 5632 16056 5684 16108
rect 9128 16056 9180 16108
rect 7288 15988 7340 16040
rect 2964 15963 3016 15972
rect 2964 15929 2973 15963
rect 2973 15929 3007 15963
rect 3007 15929 3016 15963
rect 2964 15920 3016 15929
rect 4252 15920 4304 15972
rect 9496 16192 9548 16244
rect 12808 16192 12860 16244
rect 12900 16235 12952 16244
rect 12900 16201 12909 16235
rect 12909 16201 12943 16235
rect 12943 16201 12952 16235
rect 12900 16192 12952 16201
rect 9864 16124 9916 16176
rect 14832 16192 14884 16244
rect 16764 16124 16816 16176
rect 11152 16056 11204 16108
rect 12624 16031 12676 16040
rect 12624 15997 12633 16031
rect 12633 15997 12667 16031
rect 12667 15997 12676 16031
rect 12624 15988 12676 15997
rect 15016 16099 15068 16108
rect 15016 16065 15025 16099
rect 15025 16065 15059 16099
rect 15059 16065 15068 16099
rect 15016 16056 15068 16065
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 12992 16031 13044 16040
rect 12992 15997 13001 16031
rect 13001 15997 13035 16031
rect 13035 15997 13044 16031
rect 12992 15988 13044 15997
rect 13084 16031 13136 16040
rect 13084 15997 13093 16031
rect 13093 15997 13127 16031
rect 13127 15997 13136 16031
rect 13084 15988 13136 15997
rect 14096 15988 14148 16040
rect 12808 15920 12860 15972
rect 6828 15852 6880 15904
rect 7472 15895 7524 15904
rect 7472 15861 7481 15895
rect 7481 15861 7515 15895
rect 7515 15861 7524 15895
rect 7472 15852 7524 15861
rect 8024 15852 8076 15904
rect 12532 15852 12584 15904
rect 13084 15852 13136 15904
rect 14004 15852 14056 15904
rect 16580 16056 16632 16108
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 17500 15988 17552 16040
rect 18144 15920 18196 15972
rect 15108 15852 15160 15904
rect 15752 15852 15804 15904
rect 16580 15852 16632 15904
rect 17408 15852 17460 15904
rect 18052 15852 18104 15904
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 16950 15750 17002 15802
rect 17014 15750 17066 15802
rect 17078 15750 17130 15802
rect 17142 15750 17194 15802
rect 17206 15750 17258 15802
rect 8760 15648 8812 15700
rect 9588 15648 9640 15700
rect 10140 15580 10192 15632
rect 11980 15648 12032 15700
rect 13176 15648 13228 15700
rect 4528 15555 4580 15564
rect 4528 15521 4537 15555
rect 4537 15521 4571 15555
rect 4571 15521 4580 15555
rect 4528 15512 4580 15521
rect 4988 15512 5040 15564
rect 6460 15512 6512 15564
rect 10600 15512 10652 15564
rect 11428 15512 11480 15564
rect 11704 15512 11756 15564
rect 12256 15580 12308 15632
rect 12440 15623 12492 15632
rect 12440 15589 12449 15623
rect 12449 15589 12483 15623
rect 12483 15589 12492 15623
rect 16856 15648 16908 15700
rect 12440 15580 12492 15589
rect 12164 15512 12216 15564
rect 5356 15444 5408 15496
rect 12256 15444 12308 15496
rect 13912 15487 13964 15496
rect 13912 15453 13921 15487
rect 13921 15453 13955 15487
rect 13955 15453 13964 15487
rect 13912 15444 13964 15453
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 3424 15376 3476 15428
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 4988 15351 5040 15360
rect 4988 15317 5013 15351
rect 5013 15317 5040 15351
rect 4988 15308 5040 15317
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 8852 15308 8904 15360
rect 9496 15308 9548 15360
rect 11244 15376 11296 15428
rect 11152 15308 11204 15360
rect 11336 15308 11388 15360
rect 11704 15308 11756 15360
rect 12808 15308 12860 15360
rect 13728 15308 13780 15360
rect 13820 15351 13872 15360
rect 13820 15317 13829 15351
rect 13829 15317 13863 15351
rect 13863 15317 13872 15351
rect 13820 15308 13872 15317
rect 14372 15419 14424 15428
rect 14372 15385 14381 15419
rect 14381 15385 14415 15419
rect 14415 15385 14424 15419
rect 14372 15376 14424 15385
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 17610 15206 17662 15258
rect 17674 15206 17726 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 10968 15104 11020 15156
rect 6552 15036 6604 15088
rect 10692 15036 10744 15088
rect 11152 15104 11204 15156
rect 11520 15104 11572 15156
rect 11888 15147 11940 15156
rect 11888 15113 11897 15147
rect 11897 15113 11931 15147
rect 11931 15113 11940 15147
rect 11888 15104 11940 15113
rect 11980 15147 12032 15156
rect 11980 15113 11989 15147
rect 11989 15113 12023 15147
rect 12023 15113 12032 15147
rect 11980 15104 12032 15113
rect 12072 15104 12124 15156
rect 6092 14968 6144 15020
rect 11152 15011 11204 15020
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 11612 15036 11664 15088
rect 11428 14968 11480 15020
rect 12348 15011 12400 15020
rect 12348 14977 12357 15011
rect 12357 14977 12391 15011
rect 12391 14977 12400 15011
rect 12348 14968 12400 14977
rect 14740 15011 14792 15020
rect 14740 14977 14749 15011
rect 14749 14977 14783 15011
rect 14783 14977 14792 15011
rect 14740 14968 14792 14977
rect 9588 14900 9640 14952
rect 10784 14900 10836 14952
rect 6276 14832 6328 14884
rect 5080 14764 5132 14816
rect 12072 14764 12124 14816
rect 12992 14900 13044 14952
rect 13084 14900 13136 14952
rect 16304 15036 16356 15088
rect 15384 14968 15436 15020
rect 13912 14832 13964 14884
rect 15108 14832 15160 14884
rect 16948 14832 17000 14884
rect 18696 14900 18748 14952
rect 13084 14764 13136 14816
rect 13360 14764 13412 14816
rect 15292 14807 15344 14816
rect 15292 14773 15301 14807
rect 15301 14773 15335 14807
rect 15335 14773 15344 14807
rect 15292 14764 15344 14773
rect 16764 14764 16816 14816
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 16950 14662 17002 14714
rect 17014 14662 17066 14714
rect 17078 14662 17130 14714
rect 17142 14662 17194 14714
rect 17206 14662 17258 14714
rect 6552 14603 6604 14612
rect 6552 14569 6561 14603
rect 6561 14569 6595 14603
rect 6595 14569 6604 14603
rect 6552 14560 6604 14569
rect 8392 14560 8444 14612
rect 14740 14560 14792 14612
rect 13912 14492 13964 14544
rect 14280 14492 14332 14544
rect 11704 14424 11756 14476
rect 11980 14424 12032 14476
rect 13544 14424 13596 14476
rect 15384 14424 15436 14476
rect 16028 14424 16080 14476
rect 6092 14356 6144 14408
rect 6552 14356 6604 14408
rect 6828 14356 6880 14408
rect 9404 14356 9456 14408
rect 11428 14356 11480 14408
rect 2872 14288 2924 14340
rect 2964 14263 3016 14272
rect 2964 14229 2973 14263
rect 2973 14229 3007 14263
rect 3007 14229 3016 14263
rect 2964 14220 3016 14229
rect 3056 14263 3108 14272
rect 3056 14229 3065 14263
rect 3065 14229 3099 14263
rect 3099 14229 3108 14263
rect 3056 14220 3108 14229
rect 6184 14220 6236 14272
rect 11612 14288 11664 14340
rect 14832 14356 14884 14408
rect 14464 14288 14516 14340
rect 15200 14288 15252 14340
rect 15660 14288 15712 14340
rect 12256 14263 12308 14272
rect 12256 14229 12281 14263
rect 12281 14229 12308 14263
rect 12256 14220 12308 14229
rect 12440 14263 12492 14272
rect 12440 14229 12449 14263
rect 12449 14229 12483 14263
rect 12483 14229 12492 14263
rect 12440 14220 12492 14229
rect 15844 14220 15896 14272
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 17610 14118 17662 14170
rect 17674 14118 17726 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 3056 14016 3108 14068
rect 14832 14016 14884 14068
rect 4068 13948 4120 14000
rect 5908 13948 5960 14000
rect 6552 13948 6604 14000
rect 11152 13948 11204 14000
rect 13544 13948 13596 14000
rect 2504 13923 2556 13932
rect 2504 13889 2513 13923
rect 2513 13889 2547 13923
rect 2547 13889 2556 13923
rect 2504 13880 2556 13889
rect 6184 13880 6236 13932
rect 8576 13880 8628 13932
rect 10876 13880 10928 13932
rect 13176 13880 13228 13932
rect 15200 13880 15252 13932
rect 3516 13812 3568 13864
rect 4344 13812 4396 13864
rect 5724 13812 5776 13864
rect 6368 13812 6420 13864
rect 6552 13812 6604 13864
rect 4160 13744 4212 13796
rect 8484 13812 8536 13864
rect 11152 13812 11204 13864
rect 11428 13812 11480 13864
rect 12164 13812 12216 13864
rect 14188 13812 14240 13864
rect 16120 13812 16172 13864
rect 4896 13676 4948 13728
rect 6920 13676 6972 13728
rect 7288 13676 7340 13728
rect 9036 13676 9088 13728
rect 13084 13676 13136 13728
rect 13544 13676 13596 13728
rect 15476 13676 15528 13728
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 16950 13574 17002 13626
rect 17014 13574 17066 13626
rect 17078 13574 17130 13626
rect 17142 13574 17194 13626
rect 17206 13574 17258 13626
rect 4528 13472 4580 13524
rect 6920 13472 6972 13524
rect 7472 13472 7524 13524
rect 13268 13472 13320 13524
rect 4436 13404 4488 13456
rect 10600 13404 10652 13456
rect 10968 13404 11020 13456
rect 13084 13404 13136 13456
rect 14924 13404 14976 13456
rect 2136 13311 2188 13320
rect 2136 13277 2145 13311
rect 2145 13277 2179 13311
rect 2179 13277 2188 13311
rect 2136 13268 2188 13277
rect 2412 13311 2464 13320
rect 2412 13277 2421 13311
rect 2421 13277 2455 13311
rect 2455 13277 2464 13311
rect 2412 13268 2464 13277
rect 7472 13336 7524 13388
rect 8116 13336 8168 13388
rect 2320 13243 2372 13252
rect 2320 13209 2329 13243
rect 2329 13209 2363 13243
rect 2363 13209 2372 13243
rect 2320 13200 2372 13209
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 4528 13268 4580 13320
rect 5540 13268 5592 13320
rect 6092 13268 6144 13320
rect 7104 13268 7156 13320
rect 8944 13268 8996 13320
rect 10048 13268 10100 13320
rect 10876 13268 10928 13320
rect 13452 13268 13504 13320
rect 14004 13268 14056 13320
rect 14740 13268 14792 13320
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 3516 13200 3568 13252
rect 13820 13243 13872 13252
rect 13820 13209 13829 13243
rect 13829 13209 13863 13243
rect 13863 13209 13872 13243
rect 13820 13200 13872 13209
rect 14096 13243 14148 13252
rect 14096 13209 14105 13243
rect 14105 13209 14139 13243
rect 14139 13209 14148 13243
rect 14096 13200 14148 13209
rect 16304 13200 16356 13252
rect 6000 13132 6052 13184
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 6644 13132 6696 13184
rect 9588 13132 9640 13184
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 11888 13132 11940 13184
rect 14464 13132 14516 13184
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 17610 13030 17662 13082
rect 17674 13030 17726 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 5632 12928 5684 12980
rect 7564 12928 7616 12980
rect 10140 12928 10192 12980
rect 10968 12928 11020 12980
rect 11612 12928 11664 12980
rect 12256 12928 12308 12980
rect 13268 12928 13320 12980
rect 14924 12928 14976 12980
rect 16304 12928 16356 12980
rect 18144 12928 18196 12980
rect 18420 12928 18472 12980
rect 5540 12860 5592 12912
rect 6552 12860 6604 12912
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 6184 12792 6236 12844
rect 6644 12792 6696 12844
rect 7840 12860 7892 12912
rect 10692 12860 10744 12912
rect 7104 12724 7156 12776
rect 7564 12724 7616 12776
rect 18144 12835 18196 12844
rect 18144 12801 18153 12835
rect 18153 12801 18187 12835
rect 18187 12801 18196 12835
rect 18144 12792 18196 12801
rect 3884 12656 3936 12708
rect 4160 12656 4212 12708
rect 4896 12656 4948 12708
rect 5632 12656 5684 12708
rect 7656 12656 7708 12708
rect 9128 12724 9180 12776
rect 9220 12724 9272 12776
rect 11428 12724 11480 12776
rect 11520 12724 11572 12776
rect 11704 12724 11756 12776
rect 14188 12724 14240 12776
rect 14740 12767 14792 12776
rect 14740 12733 14749 12767
rect 14749 12733 14783 12767
rect 14783 12733 14792 12767
rect 14740 12724 14792 12733
rect 9496 12656 9548 12708
rect 16212 12724 16264 12776
rect 16580 12724 16632 12776
rect 16396 12656 16448 12708
rect 4344 12631 4396 12640
rect 4344 12597 4353 12631
rect 4353 12597 4387 12631
rect 4387 12597 4396 12631
rect 4344 12588 4396 12597
rect 4712 12588 4764 12640
rect 7748 12588 7800 12640
rect 14372 12588 14424 12640
rect 15108 12588 15160 12640
rect 16764 12588 16816 12640
rect 16856 12588 16908 12640
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 16950 12486 17002 12538
rect 17014 12486 17066 12538
rect 17078 12486 17130 12538
rect 17142 12486 17194 12538
rect 17206 12486 17258 12538
rect 3884 12384 3936 12436
rect 4344 12384 4396 12436
rect 4252 12316 4304 12368
rect 4896 12316 4948 12368
rect 8392 12316 8444 12368
rect 8944 12427 8996 12436
rect 8944 12393 8953 12427
rect 8953 12393 8987 12427
rect 8987 12393 8996 12427
rect 8944 12384 8996 12393
rect 10048 12384 10100 12436
rect 10600 12384 10652 12436
rect 11704 12384 11756 12436
rect 16580 12384 16632 12436
rect 16764 12384 16816 12436
rect 3056 12248 3108 12300
rect 5264 12248 5316 12300
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 6368 12291 6420 12300
rect 6368 12257 6377 12291
rect 6377 12257 6411 12291
rect 6411 12257 6420 12291
rect 6368 12248 6420 12257
rect 6552 12291 6604 12300
rect 6552 12257 6561 12291
rect 6561 12257 6595 12291
rect 6595 12257 6604 12291
rect 6552 12248 6604 12257
rect 8300 12248 8352 12300
rect 10876 12359 10928 12368
rect 10876 12325 10885 12359
rect 10885 12325 10919 12359
rect 10919 12325 10928 12359
rect 10876 12316 10928 12325
rect 9588 12291 9640 12300
rect 9588 12257 9597 12291
rect 9597 12257 9631 12291
rect 9631 12257 9640 12291
rect 9588 12248 9640 12257
rect 2872 12180 2924 12232
rect 2504 12044 2556 12096
rect 4068 12180 4120 12232
rect 6644 12180 6696 12232
rect 6920 12180 6972 12232
rect 9036 12180 9088 12232
rect 9680 12180 9732 12232
rect 9864 12180 9916 12232
rect 14280 12316 14332 12368
rect 16304 12316 16356 12368
rect 17316 12316 17368 12368
rect 13728 12248 13780 12300
rect 14556 12248 14608 12300
rect 7104 12112 7156 12164
rect 8024 12112 8076 12164
rect 8484 12112 8536 12164
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 10416 12112 10468 12164
rect 11796 12112 11848 12164
rect 13452 12112 13504 12164
rect 13728 12112 13780 12164
rect 5080 12044 5132 12096
rect 6092 12087 6144 12096
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 6920 12044 6972 12096
rect 9588 12044 9640 12096
rect 10232 12044 10284 12096
rect 10692 12087 10744 12096
rect 10692 12053 10710 12087
rect 10710 12053 10744 12087
rect 10692 12044 10744 12053
rect 11336 12044 11388 12096
rect 11520 12044 11572 12096
rect 11888 12044 11940 12096
rect 15844 12044 15896 12096
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 17610 11942 17662 11994
rect 17674 11942 17726 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 3332 11840 3384 11892
rect 3884 11840 3936 11892
rect 6736 11840 6788 11892
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 5172 11772 5224 11824
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 2504 11704 2556 11756
rect 1860 11568 1912 11620
rect 3056 11704 3108 11756
rect 3332 11704 3384 11756
rect 4620 11704 4672 11756
rect 9680 11840 9732 11892
rect 10416 11840 10468 11892
rect 11796 11840 11848 11892
rect 13452 11840 13504 11892
rect 14096 11840 14148 11892
rect 9036 11772 9088 11824
rect 13176 11772 13228 11824
rect 8116 11704 8168 11756
rect 10416 11747 10468 11756
rect 10416 11713 10421 11747
rect 10421 11713 10455 11747
rect 10455 11713 10468 11747
rect 10416 11704 10468 11713
rect 2964 11636 3016 11688
rect 4896 11636 4948 11688
rect 6368 11636 6420 11688
rect 6552 11679 6604 11688
rect 6552 11645 6561 11679
rect 6561 11645 6595 11679
rect 6595 11645 6604 11679
rect 6552 11636 6604 11645
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 4252 11568 4304 11620
rect 6368 11500 6420 11552
rect 8668 11636 8720 11688
rect 10600 11679 10652 11688
rect 10600 11645 10609 11679
rect 10609 11645 10643 11679
rect 10643 11645 10652 11679
rect 10600 11636 10652 11645
rect 11888 11704 11940 11756
rect 11796 11636 11848 11688
rect 15568 11704 15620 11756
rect 7472 11611 7524 11620
rect 7472 11577 7481 11611
rect 7481 11577 7515 11611
rect 7515 11577 7524 11611
rect 7472 11568 7524 11577
rect 7656 11568 7708 11620
rect 9956 11568 10008 11620
rect 7104 11543 7156 11552
rect 7104 11509 7113 11543
rect 7113 11509 7147 11543
rect 7147 11509 7156 11543
rect 7104 11500 7156 11509
rect 8668 11500 8720 11552
rect 10324 11500 10376 11552
rect 11704 11500 11756 11552
rect 12992 11500 13044 11552
rect 14096 11500 14148 11552
rect 14740 11500 14792 11552
rect 17224 11500 17276 11552
rect 18144 11500 18196 11552
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 16950 11398 17002 11450
rect 17014 11398 17066 11450
rect 17078 11398 17130 11450
rect 17142 11398 17194 11450
rect 17206 11398 17258 11450
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 4528 11339 4580 11348
rect 4528 11305 4537 11339
rect 4537 11305 4571 11339
rect 4571 11305 4580 11339
rect 4528 11296 4580 11305
rect 5816 11296 5868 11348
rect 8668 11296 8720 11348
rect 9128 11296 9180 11348
rect 10600 11296 10652 11348
rect 10784 11296 10836 11348
rect 11060 11296 11112 11348
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 6552 11228 6604 11280
rect 9404 11228 9456 11280
rect 5080 11160 5132 11212
rect 6460 11160 6512 11212
rect 7472 11160 7524 11212
rect 9588 11160 9640 11212
rect 9772 11160 9824 11212
rect 3884 11092 3936 11144
rect 4160 11092 4212 11144
rect 2596 10956 2648 11008
rect 3516 10956 3568 11008
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 4436 10956 4488 11008
rect 8116 11092 8168 11144
rect 8668 11092 8720 11144
rect 8760 11092 8812 11144
rect 8944 11092 8996 11144
rect 6000 10956 6052 11008
rect 7288 11024 7340 11076
rect 6644 10956 6696 11008
rect 8116 10956 8168 11008
rect 9772 11024 9824 11076
rect 10232 11228 10284 11280
rect 11704 11228 11756 11280
rect 12256 11228 12308 11280
rect 13544 11296 13596 11348
rect 15844 11271 15896 11280
rect 15844 11237 15853 11271
rect 15853 11237 15887 11271
rect 15887 11237 15896 11271
rect 15844 11228 15896 11237
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 16856 11160 16908 11212
rect 12532 11092 12584 11144
rect 14004 11092 14056 11144
rect 16948 11092 17000 11144
rect 9036 10956 9088 11008
rect 11060 11024 11112 11076
rect 12256 11024 12308 11076
rect 14924 11024 14976 11076
rect 11980 10956 12032 11008
rect 14188 10956 14240 11008
rect 14556 10956 14608 11008
rect 16396 10956 16448 11008
rect 17316 10956 17368 11008
rect 17500 10956 17552 11008
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 17610 10854 17662 10906
rect 17674 10854 17726 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 1676 10616 1728 10668
rect 5448 10752 5500 10804
rect 5540 10752 5592 10804
rect 5632 10684 5684 10736
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 5540 10616 5592 10668
rect 5908 10616 5960 10668
rect 8760 10616 8812 10668
rect 11704 10752 11756 10804
rect 11980 10752 12032 10804
rect 14188 10752 14240 10804
rect 16212 10752 16264 10804
rect 17132 10752 17184 10804
rect 17684 10752 17736 10804
rect 9588 10684 9640 10736
rect 16672 10684 16724 10736
rect 16856 10684 16908 10736
rect 17224 10727 17276 10736
rect 17224 10693 17233 10727
rect 17233 10693 17267 10727
rect 17267 10693 17276 10727
rect 17224 10684 17276 10693
rect 17500 10684 17552 10736
rect 18696 10684 18748 10736
rect 9956 10616 10008 10668
rect 2412 10480 2464 10532
rect 9404 10548 9456 10600
rect 16672 10548 16724 10600
rect 16948 10548 17000 10600
rect 17224 10548 17276 10600
rect 17592 10548 17644 10600
rect 5264 10480 5316 10532
rect 11060 10480 11112 10532
rect 11152 10480 11204 10532
rect 13176 10480 13228 10532
rect 14188 10480 14240 10532
rect 14464 10480 14516 10532
rect 15200 10523 15252 10532
rect 15200 10489 15209 10523
rect 15209 10489 15243 10523
rect 15243 10489 15252 10523
rect 15200 10480 15252 10489
rect 15568 10480 15620 10532
rect 17500 10480 17552 10532
rect 18788 10480 18840 10532
rect 11520 10412 11572 10464
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 16212 10412 16264 10464
rect 18144 10455 18196 10464
rect 18144 10421 18153 10455
rect 18153 10421 18187 10455
rect 18187 10421 18196 10455
rect 18144 10412 18196 10421
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 16950 10310 17002 10362
rect 17014 10310 17066 10362
rect 17078 10310 17130 10362
rect 17142 10310 17194 10362
rect 17206 10310 17258 10362
rect 6644 10208 6696 10260
rect 8300 10208 8352 10260
rect 6920 10140 6972 10192
rect 10876 10208 10928 10260
rect 15568 10208 15620 10260
rect 15844 10208 15896 10260
rect 13912 10140 13964 10192
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 4896 10072 4948 10124
rect 5264 10072 5316 10124
rect 7472 10115 7524 10124
rect 7472 10081 7481 10115
rect 7481 10081 7515 10115
rect 7515 10081 7524 10115
rect 7472 10072 7524 10081
rect 8208 10072 8260 10124
rect 9588 10072 9640 10124
rect 10416 10072 10468 10124
rect 14004 10072 14056 10124
rect 14096 10072 14148 10124
rect 4252 9936 4304 9988
rect 4620 9936 4672 9988
rect 4344 9911 4396 9920
rect 4344 9877 4353 9911
rect 4353 9877 4387 9911
rect 4387 9877 4396 9911
rect 4344 9868 4396 9877
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 6736 10004 6788 10056
rect 7012 10004 7064 10056
rect 5264 9979 5316 9988
rect 5264 9945 5273 9979
rect 5273 9945 5307 9979
rect 5307 9945 5316 9979
rect 5264 9936 5316 9945
rect 5724 9936 5776 9988
rect 8116 10004 8168 10056
rect 13820 10004 13872 10056
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 16856 10140 16908 10192
rect 16948 10072 17000 10124
rect 17592 10072 17644 10124
rect 17684 10004 17736 10056
rect 18052 10004 18104 10056
rect 8760 9936 8812 9988
rect 10600 9936 10652 9988
rect 11152 9936 11204 9988
rect 5080 9868 5132 9920
rect 6552 9868 6604 9920
rect 7196 9911 7248 9920
rect 7196 9877 7205 9911
rect 7205 9877 7239 9911
rect 7239 9877 7248 9911
rect 7196 9868 7248 9877
rect 7472 9868 7524 9920
rect 8024 9868 8076 9920
rect 9772 9868 9824 9920
rect 13728 9936 13780 9988
rect 16396 9936 16448 9988
rect 12256 9868 12308 9920
rect 15844 9868 15896 9920
rect 16212 9868 16264 9920
rect 18144 9979 18196 9988
rect 18144 9945 18153 9979
rect 18153 9945 18187 9979
rect 18187 9945 18196 9979
rect 18144 9936 18196 9945
rect 18236 9911 18288 9920
rect 18236 9877 18245 9911
rect 18245 9877 18279 9911
rect 18279 9877 18288 9911
rect 18236 9868 18288 9877
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 17610 9766 17662 9818
rect 17674 9766 17726 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 3884 9664 3936 9716
rect 1768 9639 1820 9648
rect 1768 9605 1777 9639
rect 1777 9605 1811 9639
rect 1811 9605 1820 9639
rect 1768 9596 1820 9605
rect 6092 9596 6144 9648
rect 9036 9664 9088 9716
rect 10416 9664 10468 9716
rect 16120 9664 16172 9716
rect 16396 9664 16448 9716
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 5172 9571 5224 9580
rect 5172 9537 5181 9571
rect 5181 9537 5215 9571
rect 5215 9537 5224 9571
rect 5172 9528 5224 9537
rect 10784 9596 10836 9648
rect 10232 9528 10284 9580
rect 14096 9596 14148 9648
rect 14372 9596 14424 9648
rect 14464 9639 14516 9648
rect 14464 9605 14473 9639
rect 14473 9605 14507 9639
rect 14507 9605 14516 9639
rect 14464 9596 14516 9605
rect 15660 9596 15712 9648
rect 10968 9528 11020 9580
rect 4988 9460 5040 9512
rect 5080 9324 5132 9376
rect 7472 9460 7524 9512
rect 7748 9460 7800 9512
rect 8852 9503 8904 9512
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 12440 9528 12492 9580
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 14832 9528 14884 9580
rect 12348 9460 12400 9512
rect 8300 9324 8352 9376
rect 9864 9324 9916 9376
rect 10876 9324 10928 9376
rect 11244 9324 11296 9376
rect 13820 9324 13872 9376
rect 15476 9324 15528 9376
rect 15844 9324 15896 9376
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 16950 9222 17002 9274
rect 17014 9222 17066 9274
rect 17078 9222 17130 9274
rect 17142 9222 17194 9274
rect 17206 9222 17258 9274
rect 3424 9120 3476 9172
rect 3516 9052 3568 9104
rect 7380 9120 7432 9172
rect 7840 9052 7892 9104
rect 5080 8984 5132 9036
rect 6460 8984 6512 9036
rect 7012 8984 7064 9036
rect 7932 8984 7984 9036
rect 8392 9052 8444 9104
rect 9588 9052 9640 9104
rect 11060 9052 11112 9104
rect 11520 9052 11572 9104
rect 2964 8916 3016 8968
rect 3976 8916 4028 8968
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 4988 8848 5040 8900
rect 6092 8848 6144 8900
rect 7288 8916 7340 8968
rect 13728 8984 13780 9036
rect 8668 8916 8720 8968
rect 9588 8916 9640 8968
rect 11796 8916 11848 8968
rect 8760 8848 8812 8900
rect 9036 8848 9088 8900
rect 9312 8891 9364 8900
rect 9312 8857 9321 8891
rect 9321 8857 9355 8891
rect 9355 8857 9364 8891
rect 9312 8848 9364 8857
rect 11060 8848 11112 8900
rect 13084 8848 13136 8900
rect 940 8780 992 8832
rect 8392 8780 8444 8832
rect 8484 8780 8536 8832
rect 9404 8780 9456 8832
rect 10324 8780 10376 8832
rect 12532 8780 12584 8832
rect 18236 8916 18288 8968
rect 15844 8848 15896 8900
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 17610 8678 17662 8730
rect 17674 8678 17726 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 3792 8619 3844 8628
rect 3792 8585 3801 8619
rect 3801 8585 3835 8619
rect 3835 8585 3844 8619
rect 3792 8576 3844 8585
rect 5448 8576 5500 8628
rect 11152 8576 11204 8628
rect 8208 8508 8260 8560
rect 8576 8508 8628 8560
rect 3240 8440 3292 8492
rect 3976 8440 4028 8492
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 11520 8508 11572 8560
rect 14004 8508 14056 8560
rect 15936 8508 15988 8560
rect 4896 8372 4948 8424
rect 6460 8372 6512 8424
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 7380 8415 7432 8424
rect 5908 8304 5960 8356
rect 6092 8236 6144 8288
rect 7380 8381 7414 8415
rect 7414 8381 7432 8415
rect 7380 8372 7432 8381
rect 8116 8372 8168 8424
rect 13820 8372 13872 8424
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 8208 8347 8260 8356
rect 8208 8313 8217 8347
rect 8217 8313 8251 8347
rect 8251 8313 8260 8347
rect 8208 8304 8260 8313
rect 8392 8236 8444 8288
rect 8760 8236 8812 8288
rect 8852 8236 8904 8288
rect 12348 8304 12400 8356
rect 15108 8304 15160 8356
rect 18144 8347 18196 8356
rect 18144 8313 18153 8347
rect 18153 8313 18187 8347
rect 18187 8313 18196 8347
rect 18144 8304 18196 8313
rect 14832 8236 14884 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 16950 8134 17002 8186
rect 17014 8134 17066 8186
rect 17078 8134 17130 8186
rect 17142 8134 17194 8186
rect 17206 8134 17258 8186
rect 5264 8032 5316 8084
rect 6736 8032 6788 8084
rect 7012 8032 7064 8084
rect 15292 8032 15344 8084
rect 9772 7964 9824 8016
rect 16304 7964 16356 8016
rect 2412 7828 2464 7880
rect 6552 7828 6604 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 8760 7896 8812 7948
rect 12440 7896 12492 7948
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 9772 7803 9824 7812
rect 9772 7769 9781 7803
rect 9781 7769 9815 7803
rect 9815 7769 9824 7803
rect 9772 7760 9824 7769
rect 17316 7760 17368 7812
rect 5540 7692 5592 7744
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 17610 7590 17662 7642
rect 17674 7590 17726 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 3148 7488 3200 7540
rect 5356 7352 5408 7404
rect 5724 7352 5776 7404
rect 5816 7352 5868 7404
rect 7380 7420 7432 7472
rect 3976 7216 4028 7268
rect 5724 7216 5776 7268
rect 4528 7148 4580 7200
rect 6920 7352 6972 7404
rect 8024 7352 8076 7404
rect 15016 7420 15068 7472
rect 11152 7352 11204 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 13452 7352 13504 7404
rect 17408 7352 17460 7404
rect 6552 7327 6604 7336
rect 6552 7293 6561 7327
rect 6561 7293 6595 7327
rect 6595 7293 6604 7327
rect 6552 7284 6604 7293
rect 6644 7327 6696 7336
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 6644 7284 6696 7293
rect 6736 7327 6788 7336
rect 6736 7293 6745 7327
rect 6745 7293 6779 7327
rect 6779 7293 6788 7327
rect 6736 7284 6788 7293
rect 16856 7284 16908 7336
rect 7012 7216 7064 7268
rect 7104 7216 7156 7268
rect 12992 7216 13044 7268
rect 7564 7148 7616 7200
rect 8024 7148 8076 7200
rect 8300 7148 8352 7200
rect 10876 7148 10928 7200
rect 16580 7148 16632 7200
rect 17316 7148 17368 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 16950 7046 17002 7098
rect 17014 7046 17066 7098
rect 17078 7046 17130 7098
rect 17142 7046 17194 7098
rect 17206 7046 17258 7098
rect 3332 6944 3384 6996
rect 5816 6944 5868 6996
rect 5356 6876 5408 6928
rect 10048 6944 10100 6996
rect 11428 6944 11480 6996
rect 11888 6944 11940 6996
rect 12348 6944 12400 6996
rect 13728 6944 13780 6996
rect 6000 6876 6052 6928
rect 8760 6876 8812 6928
rect 12440 6876 12492 6928
rect 13452 6876 13504 6928
rect 3608 6808 3660 6860
rect 4252 6808 4304 6860
rect 4620 6740 4672 6792
rect 5816 6740 5868 6792
rect 7564 6808 7616 6860
rect 12992 6808 13044 6860
rect 16396 6808 16448 6860
rect 10416 6740 10468 6792
rect 12348 6740 12400 6792
rect 15844 6740 15896 6792
rect 3792 6672 3844 6724
rect 6736 6672 6788 6724
rect 8668 6672 8720 6724
rect 14280 6672 14332 6724
rect 14648 6672 14700 6724
rect 16764 6672 16816 6724
rect 5816 6604 5868 6656
rect 7656 6604 7708 6656
rect 13636 6604 13688 6656
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 17610 6502 17662 6554
rect 17674 6502 17726 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 2412 6332 2464 6384
rect 2872 6332 2924 6384
rect 3056 6332 3108 6384
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 1492 6264 1544 6273
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 2412 6196 2464 6248
rect 3148 6264 3200 6316
rect 6092 6400 6144 6452
rect 6184 6443 6236 6452
rect 6184 6409 6193 6443
rect 6193 6409 6227 6443
rect 6227 6409 6236 6443
rect 6184 6400 6236 6409
rect 8024 6400 8076 6452
rect 10692 6400 10744 6452
rect 3608 6332 3660 6384
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3608 6196 3660 6248
rect 940 6060 992 6112
rect 2872 6060 2924 6112
rect 4620 6332 4672 6384
rect 4712 6375 4764 6384
rect 4712 6341 4721 6375
rect 4721 6341 4755 6375
rect 4755 6341 4764 6375
rect 4712 6332 4764 6341
rect 6828 6332 6880 6384
rect 4252 6264 4304 6316
rect 6000 6264 6052 6316
rect 6184 6264 6236 6316
rect 11612 6332 11664 6384
rect 6644 6239 6696 6248
rect 6644 6205 6653 6239
rect 6653 6205 6687 6239
rect 6687 6205 6696 6239
rect 6644 6196 6696 6205
rect 6000 6128 6052 6180
rect 9128 6264 9180 6316
rect 15200 6332 15252 6384
rect 14464 6264 14516 6316
rect 18052 6264 18104 6316
rect 10140 6196 10192 6248
rect 10600 6196 10652 6248
rect 13084 6196 13136 6248
rect 13636 6196 13688 6248
rect 3792 6060 3844 6112
rect 7472 6060 7524 6112
rect 11888 6128 11940 6180
rect 12624 6128 12676 6180
rect 16028 6196 16080 6248
rect 18420 6171 18472 6180
rect 18420 6137 18429 6171
rect 18429 6137 18463 6171
rect 18463 6137 18472 6171
rect 18420 6128 18472 6137
rect 8300 6060 8352 6112
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 9404 6060 9456 6112
rect 11520 6060 11572 6112
rect 13636 6060 13688 6112
rect 14556 6060 14608 6112
rect 15108 6060 15160 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 16950 5958 17002 6010
rect 17014 5958 17066 6010
rect 17078 5958 17130 6010
rect 17142 5958 17194 6010
rect 17206 5958 17258 6010
rect 3884 5856 3936 5908
rect 3608 5788 3660 5840
rect 4528 5720 4580 5772
rect 7288 5856 7340 5908
rect 9128 5856 9180 5908
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 11336 5856 11388 5908
rect 8024 5831 8076 5840
rect 5724 5763 5776 5772
rect 5724 5729 5733 5763
rect 5733 5729 5767 5763
rect 5767 5729 5776 5763
rect 5724 5720 5776 5729
rect 6184 5720 6236 5772
rect 8024 5797 8033 5831
rect 8033 5797 8067 5831
rect 8067 5797 8076 5831
rect 8024 5788 8076 5797
rect 8116 5788 8168 5840
rect 9404 5788 9456 5840
rect 1492 5516 1544 5568
rect 4252 5584 4304 5636
rect 6828 5652 6880 5704
rect 7380 5652 7432 5704
rect 6000 5584 6052 5636
rect 7288 5584 7340 5636
rect 7564 5584 7616 5636
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 9036 5720 9088 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 9312 5652 9364 5704
rect 14924 5788 14976 5840
rect 11980 5763 12032 5772
rect 11980 5729 11989 5763
rect 11989 5729 12023 5763
rect 12023 5729 12032 5763
rect 11980 5720 12032 5729
rect 8944 5584 8996 5636
rect 11888 5584 11940 5636
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 12624 5652 12676 5704
rect 18144 5652 18196 5704
rect 14004 5584 14056 5636
rect 18420 5584 18472 5636
rect 8116 5516 8168 5568
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 8760 5516 8812 5568
rect 9220 5516 9272 5568
rect 16856 5516 16908 5568
rect 18052 5516 18104 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 17610 5414 17662 5466
rect 17674 5414 17726 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 10048 5312 10100 5364
rect 10876 5312 10928 5364
rect 14188 5312 14240 5364
rect 15016 5312 15068 5364
rect 3884 5244 3936 5296
rect 3976 5287 4028 5296
rect 3976 5253 3985 5287
rect 3985 5253 4019 5287
rect 4019 5253 4028 5287
rect 3976 5244 4028 5253
rect 5448 5244 5500 5296
rect 6368 5244 6420 5296
rect 6828 5244 6880 5296
rect 7656 5287 7708 5296
rect 3148 5176 3200 5228
rect 3608 5176 3660 5228
rect 6552 5176 6604 5228
rect 7656 5253 7665 5287
rect 7665 5253 7699 5287
rect 7699 5253 7708 5287
rect 7656 5244 7708 5253
rect 9772 5244 9824 5296
rect 11612 5244 11664 5296
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 1400 5015 1452 5024
rect 1400 4981 1409 5015
rect 1409 4981 1443 5015
rect 1443 4981 1452 5015
rect 1400 4972 1452 4981
rect 1676 4972 1728 5024
rect 3976 5108 4028 5160
rect 6276 5108 6328 5160
rect 6368 5108 6420 5160
rect 8116 5176 8168 5228
rect 9588 5176 9640 5228
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 12348 5176 12400 5228
rect 18328 5244 18380 5296
rect 8484 5108 8536 5160
rect 9772 5108 9824 5160
rect 9956 5108 10008 5160
rect 10140 5108 10192 5160
rect 12072 5108 12124 5160
rect 7288 5083 7340 5092
rect 7288 5049 7297 5083
rect 7297 5049 7331 5083
rect 7331 5049 7340 5083
rect 7288 5040 7340 5049
rect 10968 5040 11020 5092
rect 15200 5040 15252 5092
rect 5448 4972 5500 5024
rect 10232 4972 10284 5024
rect 11704 4972 11756 5024
rect 17408 4972 17460 5024
rect 17868 4972 17920 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 16950 4870 17002 4922
rect 17014 4870 17066 4922
rect 17078 4870 17130 4922
rect 17142 4870 17194 4922
rect 17206 4870 17258 4922
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 5264 4811 5316 4820
rect 5264 4777 5273 4811
rect 5273 4777 5307 4811
rect 5307 4777 5316 4811
rect 5264 4768 5316 4777
rect 7656 4768 7708 4820
rect 9496 4768 9548 4820
rect 3608 4700 3660 4752
rect 7288 4700 7340 4752
rect 16856 4768 16908 4820
rect 17408 4768 17460 4820
rect 1676 4675 1728 4684
rect 1676 4641 1685 4675
rect 1685 4641 1719 4675
rect 1719 4641 1728 4675
rect 1676 4632 1728 4641
rect 4988 4632 5040 4684
rect 5908 4632 5960 4684
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 6644 4564 6696 4616
rect 6920 4564 6972 4616
rect 7196 4564 7248 4616
rect 7472 4632 7524 4684
rect 9680 4632 9732 4684
rect 10416 4700 10468 4752
rect 3056 4496 3108 4548
rect 3424 4496 3476 4548
rect 2044 4428 2096 4480
rect 4528 4496 4580 4548
rect 5356 4496 5408 4548
rect 6828 4496 6880 4548
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 11888 4675 11940 4684
rect 11888 4641 11897 4675
rect 11897 4641 11931 4675
rect 11931 4641 11940 4675
rect 11888 4632 11940 4641
rect 11980 4632 12032 4684
rect 9956 4607 10008 4616
rect 9956 4573 9966 4607
rect 9966 4573 10000 4607
rect 10000 4573 10008 4607
rect 9956 4564 10008 4573
rect 11428 4564 11480 4616
rect 13820 4632 13872 4684
rect 15200 4607 15252 4616
rect 4436 4428 4488 4480
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 10324 4496 10376 4548
rect 15200 4573 15209 4607
rect 15209 4573 15243 4607
rect 15243 4573 15252 4607
rect 15200 4564 15252 4573
rect 11796 4496 11848 4548
rect 11980 4496 12032 4548
rect 12532 4496 12584 4548
rect 15752 4496 15804 4548
rect 8024 4428 8076 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 17610 4326 17662 4378
rect 17674 4326 17726 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 3332 4224 3384 4276
rect 2136 4199 2188 4208
rect 2136 4165 2145 4199
rect 2145 4165 2179 4199
rect 2179 4165 2188 4199
rect 2136 4156 2188 4165
rect 4804 4156 4856 4208
rect 1584 4088 1636 4140
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 2228 4088 2280 4140
rect 3608 4088 3660 4140
rect 8484 4224 8536 4276
rect 14188 4224 14240 4276
rect 17500 4224 17552 4276
rect 18420 4267 18472 4276
rect 18420 4233 18429 4267
rect 18429 4233 18463 4267
rect 18463 4233 18472 4267
rect 18420 4224 18472 4233
rect 3884 4020 3936 4072
rect 2044 3952 2096 4004
rect 2504 3995 2556 4004
rect 2504 3961 2513 3995
rect 2513 3961 2547 3995
rect 2547 3961 2556 3995
rect 2504 3952 2556 3961
rect 8392 4156 8444 4208
rect 13268 4156 13320 4208
rect 14556 4156 14608 4208
rect 18052 4199 18104 4208
rect 18052 4165 18061 4199
rect 18061 4165 18095 4199
rect 18095 4165 18104 4199
rect 18052 4156 18104 4165
rect 9956 4088 10008 4140
rect 8484 4020 8536 4072
rect 8944 4020 8996 4072
rect 11428 4020 11480 4072
rect 11796 4063 11848 4072
rect 11796 4029 11805 4063
rect 11805 4029 11839 4063
rect 11839 4029 11848 4063
rect 11796 4020 11848 4029
rect 11888 4020 11940 4072
rect 14188 4020 14240 4072
rect 15660 3952 15712 4004
rect 17592 4020 17644 4072
rect 18696 4020 18748 4072
rect 18144 3952 18196 4004
rect 3056 3884 3108 3936
rect 4344 3884 4396 3936
rect 5080 3884 5132 3936
rect 9588 3884 9640 3936
rect 9680 3884 9732 3936
rect 15292 3884 15344 3936
rect 18604 3884 18656 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 16950 3782 17002 3834
rect 17014 3782 17066 3834
rect 17078 3782 17130 3834
rect 17142 3782 17194 3834
rect 17206 3782 17258 3834
rect 1860 3680 1912 3732
rect 5540 3680 5592 3732
rect 6460 3680 6512 3732
rect 9680 3680 9732 3732
rect 11060 3680 11112 3732
rect 3700 3612 3752 3664
rect 4252 3612 4304 3664
rect 2320 3544 2372 3596
rect 4344 3544 4396 3596
rect 4896 3612 4948 3664
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 5816 3655 5868 3664
rect 5816 3621 5825 3655
rect 5825 3621 5859 3655
rect 5859 3621 5868 3655
rect 5816 3612 5868 3621
rect 11152 3655 11204 3664
rect 11152 3621 11161 3655
rect 11161 3621 11195 3655
rect 11195 3621 11204 3655
rect 11152 3612 11204 3621
rect 11336 3612 11388 3664
rect 7380 3544 7432 3596
rect 9312 3544 9364 3596
rect 11704 3544 11756 3596
rect 14556 3612 14608 3664
rect 17500 3723 17552 3732
rect 17500 3689 17509 3723
rect 17509 3689 17543 3723
rect 17543 3689 17552 3723
rect 17500 3680 17552 3689
rect 18144 3680 18196 3732
rect 12164 3544 12216 3596
rect 15108 3587 15160 3596
rect 15108 3553 15117 3587
rect 15117 3553 15151 3587
rect 15151 3553 15160 3587
rect 15108 3544 15160 3553
rect 15200 3544 15252 3596
rect 18604 3612 18656 3664
rect 18512 3544 18564 3596
rect 3884 3451 3936 3460
rect 3884 3417 3893 3451
rect 3893 3417 3927 3451
rect 3927 3417 3936 3451
rect 7288 3476 7340 3528
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 3884 3408 3936 3417
rect 4528 3408 4580 3460
rect 8852 3408 8904 3460
rect 9128 3408 9180 3460
rect 9220 3451 9272 3460
rect 9220 3417 9229 3451
rect 9229 3417 9263 3451
rect 9263 3417 9272 3451
rect 9220 3408 9272 3417
rect 10876 3408 10928 3460
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 9496 3340 9548 3392
rect 9588 3340 9640 3392
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 12256 3519 12308 3528
rect 12256 3485 12265 3519
rect 12265 3485 12299 3519
rect 12299 3485 12308 3519
rect 12256 3476 12308 3485
rect 13176 3476 13228 3528
rect 13544 3476 13596 3528
rect 17868 3476 17920 3528
rect 12072 3408 12124 3460
rect 15660 3408 15712 3460
rect 15752 3451 15804 3460
rect 15752 3417 15761 3451
rect 15761 3417 15795 3451
rect 15795 3417 15804 3451
rect 15752 3408 15804 3417
rect 17316 3408 17368 3460
rect 18144 3451 18196 3460
rect 18144 3417 18153 3451
rect 18153 3417 18187 3451
rect 18187 3417 18196 3451
rect 18144 3408 18196 3417
rect 14648 3340 14700 3392
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 17610 3238 17662 3290
rect 17674 3238 17726 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 1860 3136 1912 3188
rect 6092 3136 6144 3188
rect 3056 3068 3108 3120
rect 4068 3068 4120 3120
rect 5448 3068 5500 3120
rect 6368 3111 6420 3120
rect 6368 3077 6377 3111
rect 6377 3077 6411 3111
rect 6411 3077 6420 3111
rect 6368 3068 6420 3077
rect 6552 3179 6604 3188
rect 6552 3145 6577 3179
rect 6577 3145 6604 3179
rect 6552 3136 6604 3145
rect 1676 3000 1728 3052
rect 4252 3000 4304 3052
rect 9588 3136 9640 3188
rect 9864 3136 9916 3188
rect 12256 3136 12308 3188
rect 13360 3136 13412 3188
rect 15384 3136 15436 3188
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 9128 3068 9180 3120
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 11060 3068 11112 3120
rect 11152 3068 11204 3120
rect 14556 3068 14608 3120
rect 14924 3068 14976 3120
rect 17592 3068 17644 3120
rect 11520 3000 11572 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 4068 2932 4120 2984
rect 11336 2932 11388 2984
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 14188 3000 14240 3052
rect 15292 3043 15344 3052
rect 15292 3009 15301 3043
rect 15301 3009 15335 3043
rect 15335 3009 15344 3043
rect 15292 3000 15344 3009
rect 16764 3000 16816 3052
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 16212 2932 16264 2984
rect 16304 2932 16356 2984
rect 940 2796 992 2848
rect 8116 2864 8168 2916
rect 9220 2864 9272 2916
rect 12992 2864 13044 2916
rect 7288 2796 7340 2848
rect 11152 2796 11204 2848
rect 11336 2796 11388 2848
rect 13912 2796 13964 2848
rect 14832 2864 14884 2916
rect 16304 2839 16356 2848
rect 16304 2805 16313 2839
rect 16313 2805 16347 2839
rect 16347 2805 16356 2839
rect 16304 2796 16356 2805
rect 17500 2864 17552 2916
rect 18788 2932 18840 2984
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 16950 2694 17002 2746
rect 17014 2694 17066 2746
rect 17078 2694 17130 2746
rect 17142 2694 17194 2746
rect 17206 2694 17258 2746
rect 5908 2592 5960 2644
rect 6184 2456 6236 2508
rect 5816 2388 5868 2440
rect 10968 2592 11020 2644
rect 13636 2592 13688 2644
rect 18328 2635 18380 2644
rect 18328 2601 18337 2635
rect 18337 2601 18371 2635
rect 18371 2601 18380 2635
rect 18328 2592 18380 2601
rect 9128 2567 9180 2576
rect 9128 2533 9137 2567
rect 9137 2533 9171 2567
rect 9171 2533 9180 2567
rect 9128 2524 9180 2533
rect 11796 2524 11848 2576
rect 16304 2524 16356 2576
rect 8944 2456 8996 2508
rect 9956 2456 10008 2508
rect 8668 2388 8720 2440
rect 20 2252 72 2304
rect 2504 2252 2556 2304
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 11336 2431 11388 2440
rect 11336 2397 11345 2431
rect 11345 2397 11379 2431
rect 11379 2397 11388 2431
rect 11336 2388 11388 2397
rect 11612 2388 11664 2440
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 17960 2388 18012 2440
rect 9496 2320 9548 2372
rect 11244 2320 11296 2372
rect 12348 2252 12400 2304
rect 14188 2252 14240 2304
rect 17408 2252 17460 2304
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 17610 2150 17662 2202
rect 17674 2150 17726 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
<< metal2 >>
rect 662 19200 718 20000
rect 3882 19200 3938 20000
rect 6458 19200 6514 20000
rect 9678 19200 9734 20000
rect 12254 19200 12310 20000
rect 15474 19200 15530 20000
rect 18050 19200 18106 20000
rect 676 17270 704 19200
rect 1582 18456 1638 18465
rect 1582 18391 1638 18400
rect 1596 17338 1624 18391
rect 3896 17898 3924 19200
rect 3896 17870 4200 17898
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 4172 17338 4200 17870
rect 6472 17338 6500 19200
rect 7610 17436 7918 17445
rect 7610 17434 7616 17436
rect 7672 17434 7696 17436
rect 7752 17434 7776 17436
rect 7832 17434 7856 17436
rect 7912 17434 7918 17436
rect 7672 17382 7674 17434
rect 7854 17382 7856 17434
rect 7610 17380 7616 17382
rect 7672 17380 7696 17382
rect 7752 17380 7776 17382
rect 7832 17380 7856 17382
rect 7912 17380 7918 17382
rect 7610 17371 7918 17380
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 664 17264 716 17270
rect 664 17206 716 17212
rect 3056 17264 3108 17270
rect 3056 17206 3108 17212
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1504 16017 1532 17138
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 1490 16008 1546 16017
rect 2976 15978 3004 17002
rect 3068 16114 3096 17206
rect 9692 17202 9720 19200
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3238 16144 3294 16153
rect 3056 16108 3108 16114
rect 3238 16079 3294 16088
rect 3332 16108 3384 16114
rect 3056 16050 3108 16056
rect 1490 15943 1546 15952
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 15065 1624 15302
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 1582 15056 1638 15065
rect 2976 15042 3004 15914
rect 1582 14991 1638 15000
rect 2884 15014 3004 15042
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 2884 14346 2912 15014
rect 3068 14940 3096 16050
rect 2976 14912 3096 14940
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2976 14278 3004 14912
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 2502 13968 2558 13977
rect 2502 13903 2504 13912
rect 2556 13903 2558 13912
rect 2504 13874 2556 13880
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2148 12889 2176 13262
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2134 12880 2190 12889
rect 1584 12844 1636 12850
rect 2134 12815 2190 12824
rect 1584 12786 1636 12792
rect 1596 12345 1624 12786
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1950 11792 2006 11801
rect 1950 11727 1952 11736
rect 2004 11727 2006 11736
rect 2226 11792 2282 11801
rect 2332 11762 2360 13194
rect 2226 11727 2282 11736
rect 2320 11756 2372 11762
rect 1952 11698 2004 11704
rect 2240 11642 2268 11727
rect 2320 11698 2372 11704
rect 1860 11620 1912 11626
rect 2240 11614 2360 11642
rect 1860 11562 1912 11568
rect 1766 11248 1822 11257
rect 1766 11183 1822 11192
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1688 9586 1716 10610
rect 1780 9654 1808 11183
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 938 8936 994 8945
rect 938 8871 994 8880
rect 952 8838 980 8871
rect 940 8832 992 8838
rect 940 8774 992 8780
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 938 6216 994 6225
rect 938 6151 994 6160
rect 952 6118 980 6151
rect 940 6112 992 6118
rect 940 6054 992 6060
rect 1504 5574 1532 6258
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 3505 1440 4966
rect 1596 4146 1624 5607
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4690 1716 4966
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1398 3496 1454 3505
rect 1398 3431 1454 3440
rect 1688 3058 1716 4082
rect 1872 3738 1900 11562
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1964 6225 1992 6258
rect 1950 6216 2006 6225
rect 1950 6151 2006 6160
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2044 5160 2096 5166
rect 2042 5128 2044 5137
rect 2096 5128 2098 5137
rect 2042 5063 2098 5072
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 2056 4010 2084 4422
rect 2136 4208 2188 4214
rect 2134 4176 2136 4185
rect 2188 4176 2190 4185
rect 2332 4162 2360 11614
rect 2424 10538 2452 13262
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 2872 12232 2924 12238
rect 2870 12200 2872 12209
rect 2924 12200 2926 12209
rect 2870 12135 2926 12144
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2516 11880 2544 12038
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 2516 11852 2636 11880
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2516 10577 2544 11698
rect 2608 11014 2636 11852
rect 2976 11694 3004 14214
rect 3068 14074 3096 14214
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3054 12336 3110 12345
rect 3054 12271 3056 12280
rect 3108 12271 3110 12280
rect 3056 12242 3108 12248
rect 3068 11762 3096 12242
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 2502 10568 2558 10577
rect 2412 10532 2464 10538
rect 2502 10503 2558 10512
rect 2412 10474 2464 10480
rect 2502 10296 2558 10305
rect 2502 10231 2558 10240
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2424 6390 2452 7822
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2424 5273 2452 6190
rect 2410 5264 2466 5273
rect 2410 5199 2466 5208
rect 2240 4146 2360 4162
rect 2134 4111 2190 4120
rect 2228 4140 2360 4146
rect 2280 4134 2360 4140
rect 2228 4082 2280 4088
rect 2044 4004 2096 4010
rect 2044 3946 2096 3952
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2332 3602 2360 4134
rect 2516 4010 2544 10231
rect 3054 10024 3110 10033
rect 3054 9959 3110 9968
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2884 6118 2912 6326
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2976 6066 3004 8910
rect 3068 6390 3096 9959
rect 3160 7546 3188 13262
rect 3252 8498 3280 16079
rect 3332 16050 3384 16056
rect 3344 11898 3372 16050
rect 3424 15428 3476 15434
rect 3424 15370 3476 15376
rect 3436 14385 3464 15370
rect 3422 14376 3478 14385
rect 3422 14311 3478 14320
rect 3436 13682 3464 14311
rect 3516 13864 3568 13870
rect 3568 13812 3740 13818
rect 3516 13806 3740 13812
rect 3528 13790 3740 13806
rect 3436 13654 3648 13682
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3528 12434 3556 13194
rect 3436 12406 3556 12434
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3344 9058 3372 11698
rect 3436 9178 3464 12406
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3528 9110 3556 10950
rect 3620 10674 3648 13654
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3516 9104 3568 9110
rect 3344 9030 3464 9058
rect 3516 9046 3568 9052
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3160 6202 3188 6258
rect 3160 6174 3280 6202
rect 2976 6038 3188 6066
rect 3054 5536 3110 5545
rect 2610 5468 2918 5477
rect 3054 5471 3110 5480
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 3068 4554 3096 5471
rect 3160 5234 3188 6038
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3160 4826 3188 5170
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 3252 4434 3280 6174
rect 3068 4406 3280 4434
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 3068 3942 3096 4406
rect 3344 4282 3372 6938
rect 3436 4554 3464 9030
rect 3528 6322 3556 9046
rect 3712 7993 3740 13790
rect 3804 11354 3832 16458
rect 4080 16153 4108 17138
rect 4540 16998 4568 17138
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4356 16726 4384 16934
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 3974 15600 4030 15609
rect 3974 15535 4030 15544
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3896 12442 3924 12650
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3896 11234 3924 11834
rect 3804 11206 3924 11234
rect 3804 8634 3832 11206
rect 3884 11144 3936 11150
rect 3882 11112 3884 11121
rect 3936 11112 3938 11121
rect 3882 11047 3938 11056
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3698 7984 3754 7993
rect 3698 7919 3754 7928
rect 3698 7304 3754 7313
rect 3698 7239 3754 7248
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3620 6390 3648 6802
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5846 3648 6190
rect 3608 5840 3660 5846
rect 3608 5782 3660 5788
rect 3606 5536 3662 5545
rect 3606 5471 3662 5480
rect 3620 5234 3648 5471
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3620 4758 3648 5170
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3424 4548 3476 4554
rect 3424 4490 3476 4496
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3620 4146 3648 4694
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1872 3194 1900 3334
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 3068 3126 3096 3878
rect 3712 3670 3740 7239
rect 3804 6905 3832 8570
rect 3790 6896 3846 6905
rect 3790 6831 3846 6840
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3804 6118 3832 6666
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3896 5914 3924 9658
rect 3988 8974 4016 15535
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4080 13841 4108 13942
rect 4066 13832 4122 13841
rect 4066 13767 4122 13776
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4172 12714 4200 13738
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 4264 12374 4292 15914
rect 4540 15570 4568 16934
rect 5368 16697 5396 17070
rect 5354 16688 5410 16697
rect 5354 16623 5410 16632
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 4344 13864 4396 13870
rect 4342 13832 4344 13841
rect 4396 13832 4398 13841
rect 4342 13767 4398 13776
rect 4540 13530 4568 15506
rect 5000 15366 5028 15506
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 4988 15360 5040 15366
rect 5172 15360 5224 15366
rect 4988 15302 5040 15308
rect 5170 15328 5172 15337
rect 5224 15328 5226 15337
rect 5170 15263 5226 15272
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 4802 14512 4858 14521
rect 4802 14447 4858 14456
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4436 13456 4488 13462
rect 4436 13398 4488 13404
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4356 12442 4384 12582
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4158 12200 4214 12209
rect 4080 11218 4108 12174
rect 4158 12135 4214 12144
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4172 11150 4200 12135
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4264 11014 4292 11562
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4356 10010 4384 12378
rect 4448 11218 4476 13398
rect 4540 13326 4568 13466
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4526 12744 4582 12753
rect 4526 12679 4582 12688
rect 4540 11354 4568 12679
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4448 10713 4476 10950
rect 4434 10704 4490 10713
rect 4434 10639 4490 10648
rect 4632 10130 4660 11698
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4252 9988 4304 9994
rect 4356 9982 4476 10010
rect 4632 9994 4660 10066
rect 4252 9930 4304 9936
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 8498 4016 8910
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3988 5302 4016 7210
rect 4264 6866 4292 9930
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4264 5642 4292 6258
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4264 5545 4292 5578
rect 4250 5536 4306 5545
rect 4250 5471 4306 5480
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3896 5148 3924 5238
rect 3976 5160 4028 5166
rect 3896 5120 3976 5148
rect 3976 5102 4028 5108
rect 4250 4720 4306 4729
rect 4250 4655 4306 4664
rect 4264 4622 4292 4655
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 3884 4072 3936 4078
rect 4356 4049 4384 9862
rect 4448 4486 4476 9982
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4540 5778 4568 7142
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4632 6390 4660 6734
rect 4724 6390 4752 12582
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 3884 4014 3936 4020
rect 4342 4040 4398 4049
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3896 3466 3924 4014
rect 4342 3975 4398 3984
rect 4344 3936 4396 3942
rect 4264 3884 4344 3890
rect 4264 3878 4396 3884
rect 4264 3862 4384 3878
rect 4264 3670 4292 3862
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 4080 2990 4108 3062
rect 4264 3058 4292 3606
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4356 3097 4384 3538
rect 4540 3466 4568 4490
rect 4816 4214 4844 14447
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4908 12714 4936 13670
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4908 12434 4936 12650
rect 4908 12406 5028 12434
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4908 11694 4936 12310
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4908 8430 4936 10066
rect 5000 10062 5028 12406
rect 5092 12102 5120 14758
rect 5170 13424 5226 13433
rect 5170 13359 5226 13368
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 5092 11218 5120 12038
rect 5184 11830 5212 13359
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5092 10985 5120 11154
rect 5078 10976 5134 10985
rect 5078 10911 5134 10920
rect 5276 10538 5304 12242
rect 5368 12209 5396 15438
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 13002 5580 13262
rect 5460 12974 5580 13002
rect 5644 12986 5672 16050
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 6104 14414 6132 14962
rect 6288 14890 6316 17138
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6472 15570 6500 17002
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6276 14884 6328 14890
rect 6276 14826 6328 14832
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5632 12980 5684 12986
rect 5354 12200 5410 12209
rect 5354 12135 5410 12144
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5262 10296 5318 10305
rect 5262 10231 5318 10240
rect 5276 10130 5304 10231
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9518 5028 9998
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5092 9382 5120 9862
rect 5170 9616 5226 9625
rect 5170 9551 5172 9560
rect 5224 9551 5226 9560
rect 5172 9522 5224 9528
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5092 9042 5120 9318
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 5000 8276 5028 8842
rect 4908 8248 5028 8276
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4908 3670 4936 8248
rect 4986 5128 5042 5137
rect 4986 5063 5042 5072
rect 5000 4690 5028 5063
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5092 3942 5120 8978
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 5184 3097 5212 9522
rect 5276 8090 5304 9930
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5368 7410 5396 12135
rect 5460 10810 5488 12974
rect 5632 12922 5684 12928
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5552 10810 5580 12854
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5644 10742 5672 12650
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5552 9674 5580 10610
rect 5736 9994 5764 13806
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5552 9646 5672 9674
rect 5538 9072 5594 9081
rect 5538 9007 5594 9016
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5262 4856 5318 4865
rect 5262 4791 5264 4800
rect 5316 4791 5318 4800
rect 5264 4762 5316 4768
rect 5368 4554 5396 6870
rect 5460 5302 5488 8570
rect 5552 7750 5580 9007
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5460 3602 5488 4966
rect 5552 3738 5580 7686
rect 5644 6089 5672 9646
rect 5722 8528 5778 8537
rect 5722 8463 5778 8472
rect 5736 7410 5764 8463
rect 5828 7410 5856 11290
rect 5920 10674 5948 13942
rect 6104 13326 6132 14350
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6196 13938 6224 14214
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6012 11676 6040 13126
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6104 11801 6132 12038
rect 6090 11792 6146 11801
rect 6090 11727 6146 11736
rect 6012 11648 6132 11676
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5736 7177 5764 7210
rect 5722 7168 5778 7177
rect 5722 7103 5778 7112
rect 5828 7002 5856 7346
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5722 6896 5778 6905
rect 5722 6831 5778 6840
rect 5630 6080 5686 6089
rect 5630 6015 5686 6024
rect 5736 5778 5764 6831
rect 5816 6792 5868 6798
rect 5814 6760 5816 6769
rect 5868 6760 5870 6769
rect 5814 6695 5870 6704
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5828 3670 5856 6598
rect 5920 4690 5948 8298
rect 6012 7721 6040 10950
rect 6104 9654 6132 11648
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 6090 9480 6146 9489
rect 6090 9415 6146 9424
rect 6104 8906 6132 9415
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 5998 7712 6054 7721
rect 5998 7647 6054 7656
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 6012 6322 6040 6870
rect 6104 6458 6132 8230
rect 6196 6458 6224 12786
rect 6288 12306 6316 14826
rect 6366 13968 6422 13977
rect 6366 13903 6422 13912
rect 6380 13870 6408 13903
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 12889 6408 13126
rect 6366 12880 6422 12889
rect 6366 12815 6422 12824
rect 6472 12322 6500 15506
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6564 14618 6592 15030
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6564 14006 6592 14350
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6564 12918 6592 13806
rect 6656 13190 6684 17138
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 6950 16892 7258 16901
rect 6950 16890 6956 16892
rect 7012 16890 7036 16892
rect 7092 16890 7116 16892
rect 7172 16890 7196 16892
rect 7252 16890 7258 16892
rect 7012 16838 7014 16890
rect 7194 16838 7196 16890
rect 6950 16836 6956 16838
rect 7012 16836 7036 16838
rect 7092 16836 7116 16838
rect 7172 16836 7196 16838
rect 7252 16836 7258 16838
rect 6950 16827 7258 16836
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6932 16182 6960 16662
rect 8312 16658 8340 17070
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 7610 16348 7918 16357
rect 7610 16346 7616 16348
rect 7672 16346 7696 16348
rect 7752 16346 7776 16348
rect 7832 16346 7856 16348
rect 7912 16346 7918 16348
rect 7672 16294 7674 16346
rect 7854 16294 7856 16346
rect 7610 16292 7616 16294
rect 7672 16292 7696 16294
rect 7752 16292 7776 16294
rect 7832 16292 7856 16294
rect 7912 16292 7918 16294
rect 7610 16283 7918 16292
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7378 16008 7434 16017
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6734 15464 6790 15473
rect 6734 15399 6790 15408
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6656 12850 6684 13126
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6472 12306 6592 12322
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6368 12300 6420 12306
rect 6472 12300 6604 12306
rect 6472 12294 6552 12300
rect 6368 12242 6420 12248
rect 6552 12242 6604 12248
rect 6380 11694 6408 12242
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6368 11688 6420 11694
rect 6552 11688 6604 11694
rect 6420 11648 6500 11676
rect 6368 11630 6420 11636
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6288 7936 6316 8910
rect 6380 8498 6408 11494
rect 6472 11218 6500 11648
rect 6550 11656 6552 11665
rect 6604 11656 6606 11665
rect 6550 11591 6606 11600
rect 6564 11286 6592 11591
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6656 11014 6684 12174
rect 6748 11898 6776 15399
rect 6840 14414 6868 15846
rect 6950 15804 7258 15813
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 7300 13954 7328 15982
rect 7378 15943 7434 15952
rect 6932 13926 7328 13954
rect 6932 13734 6960 13926
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6932 12730 6960 13466
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7116 12782 7144 13262
rect 6840 12702 6960 12730
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 6840 12434 6868 12702
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 6840 12406 6960 12434
rect 6932 12238 6960 12406
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6748 10826 6776 11630
rect 6932 11540 6960 12038
rect 7116 11558 7144 12106
rect 6472 10798 6776 10826
rect 6840 11512 6960 11540
rect 7104 11552 7156 11558
rect 6472 9042 6500 10798
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6288 7908 6408 7936
rect 6274 7576 6330 7585
rect 6274 7511 6330 7520
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6012 5642 6040 6122
rect 6196 5778 6224 6258
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 6090 5536 6146 5545
rect 6090 5471 6146 5480
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 3126 5488 3538
rect 5448 3120 5500 3126
rect 4342 3088 4398 3097
rect 4252 3052 4304 3058
rect 4342 3023 4398 3032
rect 5170 3088 5226 3097
rect 5448 3062 5500 3068
rect 5170 3023 5226 3032
rect 4252 2994 4304 3000
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 940 2848 992 2854
rect 938 2816 940 2825
rect 992 2816 994 2825
rect 938 2751 994 2760
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 5920 2650 5948 4626
rect 6104 4593 6132 5471
rect 6090 4584 6146 4593
rect 6090 4519 6146 4528
rect 6104 3194 6132 4519
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6196 2514 6224 5714
rect 6288 5166 6316 7511
rect 6380 5302 6408 7908
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 3126 6408 5102
rect 6472 3738 6500 8366
rect 6564 7886 6592 9862
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6550 7712 6606 7721
rect 6550 7647 6606 7656
rect 6564 7342 6592 7647
rect 6656 7342 6684 10202
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6748 8090 6776 9998
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7721 6776 7822
rect 6734 7712 6790 7721
rect 6734 7647 6790 7656
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6550 7032 6606 7041
rect 6550 6967 6606 6976
rect 6564 5234 6592 6967
rect 6656 6474 6684 7278
rect 6748 7177 6776 7278
rect 6734 7168 6790 7177
rect 6734 7103 6790 7112
rect 6734 6896 6790 6905
rect 6734 6831 6790 6840
rect 6748 6730 6776 6831
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6656 6446 6776 6474
rect 6642 6352 6698 6361
rect 6642 6287 6698 6296
rect 6656 6254 6684 6287
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6642 6080 6698 6089
rect 6642 6015 6698 6024
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6656 4622 6684 6015
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6748 4536 6776 6446
rect 6840 6390 6868 11512
rect 7104 11494 7156 11500
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 7300 11082 7328 13670
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6932 9489 6960 10134
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6918 9480 6974 9489
rect 6918 9415 6974 9424
rect 7024 9364 7052 9998
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9761 7236 9862
rect 7194 9752 7250 9761
rect 7194 9687 7250 9696
rect 7392 9602 7420 15943
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7484 13530 7512 15846
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7484 11626 7512 13330
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7610 13019 7918 13028
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7576 12782 7604 12922
rect 7840 12912 7892 12918
rect 7668 12872 7840 12900
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7668 12714 7696 12872
rect 7840 12854 7892 12860
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7760 12481 7788 12582
rect 7746 12472 7802 12481
rect 7746 12407 7802 12416
rect 8036 12170 8064 15846
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8666 15056 8722 15065
rect 8666 14991 8722 15000
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8206 13832 8262 13841
rect 8206 13767 8262 13776
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7610 11931 7918 11940
rect 8128 11762 8156 13330
rect 8116 11756 8168 11762
rect 8036 11716 8116 11744
rect 7654 11656 7710 11665
rect 7472 11620 7524 11626
rect 7654 11591 7656 11600
rect 7472 11562 7524 11568
rect 7708 11591 7710 11600
rect 7656 11562 7708 11568
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7484 10130 7512 11154
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 8036 9926 8064 11716
rect 8116 11698 8168 11704
rect 8114 11656 8170 11665
rect 8114 11591 8170 11600
rect 8128 11150 8156 11591
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10062 8156 10950
rect 8220 10130 8248 13767
rect 8404 12374 8432 14554
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8392 12368 8444 12374
rect 8496 12345 8524 13806
rect 8392 12310 8444 12316
rect 8482 12336 8538 12345
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8312 10266 8340 12242
rect 8404 10588 8432 12310
rect 8482 12271 8538 12280
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 10713 8524 12106
rect 8482 10704 8538 10713
rect 8482 10639 8538 10648
rect 8404 10560 8524 10588
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8298 9888 8354 9897
rect 7484 9704 7512 9862
rect 7610 9820 7918 9829
rect 8298 9823 8354 9832
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 8312 9704 8340 9823
rect 7484 9676 7880 9704
rect 7392 9574 7788 9602
rect 7760 9518 7788 9574
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7024 9336 7328 9364
rect 7484 9353 7512 9454
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 7300 9160 7328 9336
rect 7470 9344 7526 9353
rect 7470 9279 7526 9288
rect 7470 9208 7526 9217
rect 7208 9132 7328 9160
rect 7380 9172 7432 9178
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7024 8430 7052 8978
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 7208 8276 7236 9132
rect 7470 9143 7526 9152
rect 7380 9114 7432 9120
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7300 8498 7328 8910
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7392 8430 7420 9114
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7208 8248 7328 8276
rect 7300 8242 7328 8248
rect 7300 8214 7420 8242
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6918 7576 6974 7585
rect 6918 7511 6974 7520
rect 6932 7410 6960 7511
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7024 7274 7052 8026
rect 7102 7848 7158 7857
rect 7102 7783 7158 7792
rect 7286 7848 7342 7857
rect 7286 7783 7342 7792
rect 7116 7274 7144 7783
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 7300 5914 7328 7783
rect 7392 7478 7420 8214
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6826 5808 6882 5817
rect 6826 5743 6882 5752
rect 6840 5710 6868 5743
rect 7392 5710 7420 7414
rect 7484 7290 7512 9143
rect 7852 9110 7880 9676
rect 8220 9676 8340 9704
rect 8220 9636 8248 9676
rect 8496 9674 8524 10560
rect 8588 10033 8616 13874
rect 8680 11694 8708 14991
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11354 8708 11494
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8772 11150 8800 15642
rect 8852 15360 8904 15366
rect 9140 15337 9168 16050
rect 8852 15302 8904 15308
rect 9126 15328 9182 15337
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8760 11144 8812 11150
rect 8864 11121 8892 15302
rect 9126 15263 9182 15272
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8956 12442 8984 13262
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 9048 12238 9076 13670
rect 9232 12782 9260 16730
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9140 12434 9168 12718
rect 9140 12406 9260 12434
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9048 11830 9076 12174
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8944 11144 8996 11150
rect 8760 11086 8812 11092
rect 8850 11112 8906 11121
rect 8574 10024 8630 10033
rect 8574 9959 8630 9968
rect 8680 9761 8708 11086
rect 9140 11121 9168 11290
rect 8944 11086 8996 11092
rect 9126 11112 9182 11121
rect 8850 11047 8906 11056
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8772 9994 8800 10610
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8666 9752 8722 9761
rect 8666 9687 8722 9696
rect 7930 9616 7986 9625
rect 7930 9551 7986 9560
rect 8036 9608 8248 9636
rect 8404 9646 8524 9674
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7944 9042 7972 9551
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 8036 7410 8064 9608
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8206 8664 8262 8673
rect 8206 8599 8262 8608
rect 8220 8566 8248 8599
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7484 7262 7696 7290
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 6866 7604 7142
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7576 6644 7604 6802
rect 7668 6662 7696 7262
rect 8024 7200 8076 7206
rect 8128 7188 8156 8366
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8220 7313 8248 8298
rect 8206 7304 8262 7313
rect 8206 7239 8262 7248
rect 8312 7206 8340 9318
rect 8404 9110 8432 9646
rect 8864 9602 8892 11047
rect 8772 9574 8892 9602
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8404 8294 8432 8774
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8390 7984 8446 7993
rect 8390 7919 8446 7928
rect 8300 7200 8352 7206
rect 8128 7160 8248 7188
rect 8024 7142 8076 7148
rect 7484 6616 7604 6644
rect 7656 6656 7708 6662
rect 7484 6202 7512 6616
rect 7656 6598 7708 6604
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 8036 6458 8064 7142
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7484 6174 7604 6202
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6840 4808 6868 5238
rect 7300 5098 7328 5578
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 6840 4780 6960 4808
rect 6932 4622 6960 4780
rect 7300 4758 7328 5034
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7484 4690 7512 6054
rect 7576 5642 7604 6174
rect 7838 5944 7894 5953
rect 7838 5879 7894 5888
rect 7852 5710 7880 5879
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 7656 5296 7708 5302
rect 7654 5264 7656 5273
rect 7708 5264 7710 5273
rect 7654 5199 7710 5208
rect 7654 4856 7710 4865
rect 7654 4791 7656 4800
rect 7708 4791 7710 4800
rect 7656 4762 7708 4768
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 6828 4548 6880 4554
rect 6748 4508 6828 4536
rect 6828 4490 6880 4496
rect 7208 4298 7236 4558
rect 8036 4486 8064 5782
rect 8128 5574 8156 5782
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7208 4270 7328 4298
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 7300 3534 7328 4270
rect 7392 3602 7420 4422
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6564 2961 6592 3130
rect 6550 2952 6606 2961
rect 6550 2887 6606 2896
rect 7300 2854 7328 3470
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 8128 2922 8156 5170
rect 8220 4729 8248 7160
rect 8300 7142 8352 7148
rect 8298 6216 8354 6225
rect 8298 6151 8354 6160
rect 8312 6118 8340 6151
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8206 4720 8262 4729
rect 8206 4655 8262 4664
rect 8312 2961 8340 5510
rect 8404 4214 8432 7919
rect 8496 5166 8524 8774
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8496 4282 8524 5102
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8392 4208 8444 4214
rect 8588 4162 8616 8502
rect 8680 6730 8708 8910
rect 8772 8906 8800 9574
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8864 8294 8892 9454
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8772 8106 8800 8230
rect 8772 8078 8892 8106
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8772 6934 8800 7890
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8680 5953 8708 6666
rect 8758 6624 8814 6633
rect 8758 6559 8814 6568
rect 8772 6089 8800 6559
rect 8758 6080 8814 6089
rect 8758 6015 8814 6024
rect 8666 5944 8722 5953
rect 8666 5879 8722 5888
rect 8392 4150 8444 4156
rect 8496 4134 8616 4162
rect 8496 4078 8524 4134
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8298 2952 8354 2961
rect 8116 2916 8168 2922
rect 8298 2887 8354 2896
rect 8116 2858 8168 2864
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 8680 2446 8708 5879
rect 8772 5574 8800 6015
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8864 3466 8892 8078
rect 8956 5642 8984 11086
rect 9126 11047 9182 11056
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 9722 9076 10950
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9048 5778 9076 8842
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5914 9168 6258
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 9232 5574 9260 12406
rect 9324 8906 9352 16730
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9508 15366 9536 16186
rect 9876 16182 9904 16526
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9600 14958 9628 15642
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9416 11286 9444 14350
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9416 8838 9444 10542
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 8537 9444 8774
rect 9402 8528 9458 8537
rect 9402 8463 9458 8472
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9324 5710 9352 6054
rect 9416 5846 9444 6054
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9402 5128 9458 5137
rect 9402 5063 9458 5072
rect 9310 4176 9366 4185
rect 9310 4111 9366 4120
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8956 3534 8984 4014
rect 9324 3602 9352 4111
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8956 2514 8984 3470
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9140 3126 9168 3402
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 9232 2922 9260 3402
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9128 2576 9180 2582
rect 9126 2544 9128 2553
rect 9180 2544 9182 2553
rect 8944 2508 8996 2514
rect 9126 2479 9182 2488
rect 8944 2450 8996 2456
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 32 800 60 2246
rect 2516 1170 2544 2246
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 2516 1142 2636 1170
rect 2608 800 2636 1142
rect 5828 800 5856 2382
rect 9416 2360 9444 5063
rect 9508 4826 9536 12650
rect 9600 12306 9628 13126
rect 9968 12434 9996 16934
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 13326 10088 16526
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10152 13138 10180 15574
rect 10060 13110 10180 13138
rect 10060 12442 10088 13110
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 9784 12406 9996 12434
rect 10048 12436 10100 12442
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11218 9628 12038
rect 9692 11898 9720 12174
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9692 11393 9720 11834
rect 9784 11529 9812 12406
rect 10048 12378 10100 12384
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9770 11520 9826 11529
rect 9770 11455 9826 11464
rect 9678 11384 9734 11393
rect 9678 11319 9734 11328
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9772 11212 9824 11218
rect 9876 11200 9904 12174
rect 10046 11928 10102 11937
rect 10046 11863 10102 11872
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9824 11172 9904 11200
rect 9772 11154 9824 11160
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9784 10826 9812 11018
rect 9692 10798 9812 10826
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9600 10130 9628 10678
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9600 8974 9628 9046
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9600 5234 9628 8910
rect 9692 5778 9720 10798
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9784 8022 9812 9862
rect 9876 9382 9904 11172
rect 9968 10674 9996 11562
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9862 8120 9918 8129
rect 9862 8055 9918 8064
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9784 5302 9812 7754
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9678 4720 9734 4729
rect 9678 4655 9680 4664
rect 9732 4655 9734 4664
rect 9680 4626 9732 4632
rect 9784 4622 9812 5102
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9600 3641 9628 3878
rect 9692 3738 9720 3878
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9586 3632 9642 3641
rect 9586 3567 9642 3576
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9508 3058 9536 3334
rect 9600 3194 9628 3334
rect 9876 3194 9904 8055
rect 9968 5166 9996 10610
rect 10060 7002 10088 11863
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10152 6338 10180 12922
rect 10244 12345 10272 16390
rect 10322 14240 10378 14249
rect 10322 14175 10378 14184
rect 10230 12336 10286 12345
rect 10230 12271 10286 12280
rect 10232 12096 10284 12102
rect 10336 12084 10364 14175
rect 10428 12434 10456 16934
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10612 15337 10640 15506
rect 10598 15328 10654 15337
rect 10598 15263 10654 15272
rect 10782 15192 10838 15201
rect 10782 15127 10838 15136
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10704 14793 10732 15030
rect 10796 14958 10824 15127
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10690 14784 10746 14793
rect 10690 14719 10746 14728
rect 10888 13938 10916 17274
rect 12268 17270 12296 19200
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12610 17371 12918 17380
rect 15488 17338 15516 19200
rect 17866 18456 17922 18465
rect 17866 18391 17922 18400
rect 17880 17626 17908 18391
rect 17880 17598 18000 17626
rect 17610 17436 17918 17445
rect 17610 17434 17616 17436
rect 17672 17434 17696 17436
rect 17752 17434 17776 17436
rect 17832 17434 17856 17436
rect 17912 17434 17918 17436
rect 17672 17382 17674 17434
rect 17854 17382 17856 17434
rect 17610 17380 17616 17382
rect 17672 17380 17696 17382
rect 17752 17380 17776 17382
rect 17832 17380 17856 17382
rect 17912 17380 17918 17382
rect 17610 17371 17918 17380
rect 17972 17338 18000 17598
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 11950 16892 12258 16901
rect 11950 16890 11956 16892
rect 12012 16890 12036 16892
rect 12092 16890 12116 16892
rect 12172 16890 12196 16892
rect 12252 16890 12258 16892
rect 12012 16838 12014 16890
rect 12194 16838 12196 16890
rect 11950 16836 11956 16838
rect 12012 16836 12036 16838
rect 12092 16836 12116 16838
rect 12172 16836 12196 16838
rect 12252 16836 12258 16838
rect 11950 16827 12258 16836
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10980 13462 11008 15098
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10968 13456 11020 13462
rect 10968 13398 11020 13404
rect 10612 12442 10640 13398
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12918 10732 13126
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10888 12458 10916 13262
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10600 12436 10652 12442
rect 10428 12406 10548 12434
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10284 12056 10364 12084
rect 10232 12038 10284 12044
rect 10428 11898 10456 12106
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10428 11762 10456 11834
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10324 11552 10376 11558
rect 10376 11512 10456 11540
rect 10324 11494 10376 11500
rect 10428 11393 10456 11512
rect 10414 11384 10470 11393
rect 10414 11319 10470 11328
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10244 11121 10272 11222
rect 10324 11144 10376 11150
rect 10230 11112 10286 11121
rect 10376 11104 10456 11132
rect 10324 11086 10376 11092
rect 10230 11047 10286 11056
rect 10230 10976 10286 10985
rect 10230 10911 10286 10920
rect 10244 9586 10272 10911
rect 10428 10130 10456 11104
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10428 9722 10456 10066
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10520 9489 10548 12406
rect 10600 12378 10652 12384
rect 10796 12430 10916 12458
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10612 11529 10640 11630
rect 10598 11520 10654 11529
rect 10598 11455 10654 11464
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10612 9994 10640 11290
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10506 9480 10562 9489
rect 10506 9415 10562 9424
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10152 6310 10272 6338
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10152 5914 10180 6190
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 10060 4690 10088 5306
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9956 4616 10008 4622
rect 9954 4584 9956 4593
rect 10152 4593 10180 5102
rect 10244 5030 10272 6310
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10008 4584 10010 4593
rect 9954 4519 10010 4528
rect 10138 4584 10194 4593
rect 10336 4554 10364 8774
rect 10612 8650 10640 9930
rect 10520 8622 10640 8650
rect 10520 8498 10548 8622
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10428 4758 10456 6734
rect 10612 6254 10640 8622
rect 10704 6458 10732 12038
rect 10796 11354 10824 12430
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10888 10266 10916 12310
rect 10980 11121 11008 12922
rect 11072 11506 11100 16458
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11164 15609 11192 16050
rect 11150 15600 11206 15609
rect 11150 15535 11206 15544
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11704 15564 11756 15570
rect 11808 15552 11836 16594
rect 12820 16590 12848 16934
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 13174 16552 13230 16561
rect 12992 16516 13044 16522
rect 13174 16487 13230 16496
rect 12992 16458 13044 16464
rect 12610 16348 12918 16357
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12900 16244 12952 16250
rect 13004 16232 13032 16458
rect 12952 16204 13032 16232
rect 12900 16186 12952 16192
rect 12820 16153 12848 16186
rect 12622 16144 12678 16153
rect 12622 16079 12678 16088
rect 12806 16144 12862 16153
rect 12806 16079 12862 16088
rect 12636 16046 12664 16079
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 12532 15904 12584 15910
rect 12636 15881 12664 15982
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12532 15846 12584 15852
rect 12622 15872 12678 15881
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11992 15609 12020 15642
rect 12256 15632 12308 15638
rect 11978 15600 12034 15609
rect 11808 15524 11928 15552
rect 12256 15574 12308 15580
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 11978 15535 12034 15544
rect 12164 15564 12216 15570
rect 11704 15506 11756 15512
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11164 15162 11192 15302
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11164 14006 11192 14962
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11164 11642 11192 13806
rect 11256 11744 11284 15370
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11348 12102 11376 15302
rect 11440 15026 11468 15506
rect 11716 15450 11744 15506
rect 11716 15422 11836 15450
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11428 14408 11480 14414
rect 11426 14376 11428 14385
rect 11480 14376 11482 14385
rect 11426 14311 11482 14320
rect 11440 13870 11468 14311
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11532 12782 11560 15098
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11624 14793 11652 15030
rect 11610 14784 11666 14793
rect 11610 14719 11666 14728
rect 11716 14482 11744 15302
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11612 14340 11664 14346
rect 11612 14282 11664 14288
rect 11624 12986 11652 14282
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11808 12866 11836 15422
rect 11900 15201 11928 15524
rect 11886 15192 11942 15201
rect 11992 15162 12020 15535
rect 12164 15506 12216 15512
rect 11886 15127 11888 15136
rect 11940 15127 11942 15136
rect 11980 15156 12032 15162
rect 11888 15098 11940 15104
rect 11980 15098 12032 15104
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12084 14822 12112 15098
rect 12176 15065 12204 15506
rect 12268 15502 12296 15574
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12452 15337 12480 15574
rect 12438 15328 12494 15337
rect 12438 15263 12494 15272
rect 12162 15056 12218 15065
rect 12162 14991 12218 15000
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11950 14716 12258 14725
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 11978 14512 12034 14521
rect 11978 14447 11980 14456
rect 12032 14447 12034 14456
rect 11980 14418 12032 14424
rect 12360 14362 12388 14962
rect 12176 14334 12388 14362
rect 12176 13870 12204 14334
rect 12256 14272 12308 14278
rect 12440 14272 12492 14278
rect 12308 14232 12388 14260
rect 12256 14214 12308 14220
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11624 12838 11836 12866
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11256 11716 11376 11744
rect 11164 11614 11284 11642
rect 11072 11478 11192 11506
rect 11058 11384 11114 11393
rect 11058 11319 11060 11328
rect 11112 11319 11114 11328
rect 11060 11290 11112 11296
rect 11058 11248 11114 11257
rect 11058 11183 11114 11192
rect 10966 11112 11022 11121
rect 11072 11082 11100 11183
rect 10966 11047 11022 11056
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11164 10538 11192 11478
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10138 4519 10194 4528
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9968 2514 9996 4082
rect 10796 4049 10824 9590
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 7698 10916 9318
rect 10980 7886 11008 9522
rect 11072 9110 11100 10474
rect 11256 10169 11284 11614
rect 11242 10160 11298 10169
rect 11242 10095 11298 10104
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10888 7670 11008 7698
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10888 5370 10916 7142
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10874 5128 10930 5137
rect 10980 5098 11008 7670
rect 11072 6769 11100 8842
rect 11164 8634 11192 9930
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11058 6760 11114 6769
rect 11058 6695 11114 6704
rect 11164 6610 11192 7346
rect 11072 6582 11192 6610
rect 10874 5063 10930 5072
rect 10968 5092 11020 5098
rect 10782 4040 10838 4049
rect 10782 3975 10838 3984
rect 10888 3466 10916 5063
rect 10968 5034 11020 5040
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10980 2650 11008 5034
rect 11072 3738 11100 6582
rect 11150 3768 11206 3777
rect 11060 3732 11112 3738
rect 11150 3703 11206 3712
rect 11060 3674 11112 3680
rect 11072 3126 11100 3674
rect 11164 3670 11192 3703
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11164 2854 11192 3062
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 11256 2378 11284 9318
rect 11348 5914 11376 11716
rect 11440 7002 11468 12718
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11532 10470 11560 12038
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11532 8566 11560 9046
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11624 7018 11652 12838
rect 11704 12776 11756 12782
rect 11900 12764 11928 13126
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12268 12889 12296 12922
rect 12254 12880 12310 12889
rect 12254 12815 12310 12824
rect 11704 12718 11756 12724
rect 11808 12736 11928 12764
rect 11716 12442 11744 12718
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11808 12322 11836 12736
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11950 12475 12258 12484
rect 11716 12294 11836 12322
rect 11716 11558 11744 12294
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11808 11898 11836 12106
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11900 11937 11928 12038
rect 11886 11928 11942 11937
rect 11796 11892 11848 11898
rect 11886 11863 11942 11872
rect 11796 11834 11848 11840
rect 11900 11762 11928 11863
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11286 11744 11494
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11532 6990 11652 7018
rect 11426 6488 11482 6497
rect 11426 6423 11482 6432
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11440 4865 11468 6423
rect 11532 6118 11560 6990
rect 11716 6882 11744 10746
rect 11808 8974 11836 11630
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 12256 11280 12308 11286
rect 12254 11248 12256 11257
rect 12308 11248 12310 11257
rect 12254 11183 12310 11192
rect 12268 11082 12296 11183
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11992 10810 12020 10950
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11950 10299 12258 10308
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12268 9364 12296 9862
rect 12360 9518 12388 14232
rect 12440 14214 12492 14220
rect 12452 9586 12480 14214
rect 12544 11150 12572 15846
rect 12622 15807 12678 15816
rect 12820 15366 12848 15914
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 13004 15042 13032 15982
rect 13096 15910 13124 15982
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13188 15706 13216 16487
rect 13266 15872 13322 15881
rect 13266 15807 13322 15816
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 12912 15014 13124 15042
rect 12912 14385 12940 15014
rect 13096 14958 13124 15014
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12898 14376 12954 14385
rect 12898 14311 12954 14320
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 13004 12753 13032 14894
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 13734 13124 14758
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 12990 12744 13046 12753
rect 12990 12679 13046 12688
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12610 10843 12918 10852
rect 12530 10160 12586 10169
rect 12530 10095 12586 10104
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12268 9336 12388 9364
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11624 6854 11744 6882
rect 11624 6497 11652 6854
rect 11702 6760 11758 6769
rect 11702 6695 11758 6704
rect 11610 6488 11666 6497
rect 11610 6423 11666 6432
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11426 4856 11482 4865
rect 11348 4814 11426 4842
rect 11348 3670 11376 4814
rect 11426 4791 11482 4800
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11440 4078 11468 4558
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11532 3058 11560 6054
rect 11624 5302 11652 6326
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11716 5114 11744 6695
rect 11624 5086 11744 5114
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11624 2990 11652 5086
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4162 11744 4966
rect 11808 4554 11836 8910
rect 12360 8362 12388 9336
rect 12452 8650 12480 9415
rect 12544 8838 12572 10095
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 12452 8622 12572 8650
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11950 8123 12258 8132
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12452 7410 12480 7890
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 11900 6186 11928 6938
rect 12360 6798 12388 6938
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 11888 6180 11940 6186
rect 11888 6122 11940 6128
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 12360 5896 12388 6734
rect 11992 5868 12388 5896
rect 11992 5778 12020 5868
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12164 5704 12216 5710
rect 12084 5664 12164 5692
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11900 5234 11928 5578
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 12084 5166 12112 5664
rect 12164 5646 12216 5652
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 11886 4720 11942 4729
rect 11886 4655 11888 4664
rect 11940 4655 11942 4664
rect 11980 4684 12032 4690
rect 11888 4626 11940 4632
rect 11980 4626 12032 4632
rect 11992 4554 12020 4626
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11716 4134 11928 4162
rect 11900 4078 11928 4134
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11808 3913 11836 4014
rect 11794 3904 11850 3913
rect 11794 3839 11850 3848
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 11716 3058 11744 3538
rect 11888 3528 11940 3534
rect 11886 3496 11888 3505
rect 11940 3496 11942 3505
rect 11886 3431 11942 3440
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12084 3097 12112 3402
rect 12176 3233 12204 3538
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12162 3224 12218 3233
rect 12268 3194 12296 3470
rect 12360 3233 12388 5170
rect 12346 3224 12402 3233
rect 12162 3159 12218 3168
rect 12256 3188 12308 3194
rect 12346 3159 12402 3168
rect 12452 3176 12480 6870
rect 12544 4554 12572 8622
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 13004 7274 13032 11494
rect 13096 8906 13124 13398
rect 13188 11830 13216 13874
rect 13280 13530 13308 15807
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12636 5710 12664 6122
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 12256 3130 12308 3136
rect 12070 3088 12126 3097
rect 11704 3052 11756 3058
rect 12070 3023 12126 3032
rect 11704 2994 11756 3000
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11794 2952 11850 2961
rect 11348 2854 11376 2926
rect 11794 2887 11850 2896
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11348 2446 11376 2790
rect 11808 2582 11836 2887
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 9496 2372 9548 2378
rect 9416 2332 9496 2360
rect 9496 2314 9548 2320
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 8496 1170 8524 2246
rect 8404 1142 8524 1170
rect 8404 800 8432 1142
rect 11624 800 11652 2382
rect 12360 2310 12388 3159
rect 12452 3148 12572 3176
rect 12544 3097 12572 3148
rect 12530 3088 12586 3097
rect 12530 3023 12586 3032
rect 13004 2922 13032 6802
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13096 3058 13124 6190
rect 13188 3534 13216 10474
rect 13280 4214 13308 12922
rect 13372 11665 13400 14758
rect 13556 14482 13584 16934
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13556 14006 13584 14418
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13464 12170 13492 13262
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13358 11656 13414 11665
rect 13358 11591 13414 11600
rect 13358 10704 13414 10713
rect 13358 10639 13414 10648
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13372 3194 13400 10639
rect 13464 8537 13492 11834
rect 13556 11354 13584 13670
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13648 10577 13676 16390
rect 14016 15910 14044 17138
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13820 15360 13872 15366
rect 13924 15337 13952 15438
rect 13820 15302 13872 15308
rect 13910 15328 13966 15337
rect 13740 12306 13768 15302
rect 13832 13410 13860 15302
rect 13910 15263 13966 15272
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13924 14550 13952 14826
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13832 13382 13952 13410
rect 13818 13288 13874 13297
rect 13818 13223 13820 13232
rect 13872 13223 13874 13232
rect 13820 13194 13872 13200
rect 13924 12434 13952 13382
rect 14016 13326 14044 15846
rect 14108 15502 14136 15982
rect 14292 15609 14320 16526
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14844 16153 14872 16186
rect 14830 16144 14886 16153
rect 14830 16079 14886 16088
rect 14278 15600 14334 15609
rect 14278 15535 14334 15544
rect 14096 15496 14148 15502
rect 14148 15456 14228 15484
rect 14096 15438 14148 15444
rect 14200 13870 14228 15456
rect 14370 15464 14426 15473
rect 14370 15399 14372 15408
rect 14424 15399 14426 15408
rect 14372 15370 14424 15376
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14752 14618 14780 14962
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 13832 12406 13952 12434
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13634 10568 13690 10577
rect 13634 10503 13690 10512
rect 13740 10452 13768 12106
rect 13556 10424 13768 10452
rect 13450 8528 13506 8537
rect 13450 8463 13506 8472
rect 13556 8378 13584 10424
rect 13634 10296 13690 10305
rect 13634 10231 13690 10240
rect 13464 8350 13584 8378
rect 13464 7410 13492 8350
rect 13542 8256 13598 8265
rect 13542 8191 13598 8200
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13464 6934 13492 7346
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 13556 3534 13584 8191
rect 13648 6746 13676 10231
rect 13832 10062 13860 12406
rect 14108 12322 14136 13194
rect 14200 12782 14228 13806
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14292 12374 14320 14486
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14476 13190 14504 14282
rect 14752 13326 14780 14554
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14844 14074 14872 14350
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 13924 12294 14136 12322
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 13924 10198 13952 12294
rect 14096 12232 14148 12238
rect 14094 12200 14096 12209
rect 14280 12232 14332 12238
rect 14148 12200 14150 12209
rect 14280 12174 14332 12180
rect 14094 12135 14150 12144
rect 14108 11898 14136 12135
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14004 11144 14056 11150
rect 14108 11132 14136 11494
rect 14056 11104 14136 11132
rect 14004 11086 14056 11092
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13740 9042 13768 9930
rect 13832 9382 13860 9998
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13832 8616 13860 9318
rect 13740 8588 13860 8616
rect 13740 7002 13768 8588
rect 13818 8528 13874 8537
rect 13818 8463 13874 8472
rect 13832 8430 13860 8463
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13648 6718 13768 6746
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 6254 13676 6598
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12992 2916 13044 2922
rect 12992 2858 13044 2864
rect 13648 2650 13676 6054
rect 13740 5137 13768 6718
rect 13818 6216 13874 6225
rect 13818 6151 13874 6160
rect 13726 5128 13782 5137
rect 13726 5063 13782 5072
rect 13832 4690 13860 6151
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13924 2854 13952 10134
rect 14016 10130 14044 11086
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10810 14228 10950
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14108 9654 14136 10066
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 14016 8430 14044 8502
rect 14108 8430 14136 9590
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14016 5642 14044 8366
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 14200 5370 14228 10474
rect 14292 6730 14320 12174
rect 14384 9654 14412 12582
rect 14476 10538 14504 13126
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14568 11014 14596 12242
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14476 6322 14504 9590
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14568 6118 14596 9522
rect 14660 6905 14688 13126
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14752 11558 14780 12718
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14844 9586 14872 14010
rect 14936 13462 14964 17070
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15212 16114 15240 17002
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15028 15337 15056 16050
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15014 15328 15070 15337
rect 15014 15263 15070 15272
rect 15120 14890 15148 15846
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 14924 13456 14976 13462
rect 14924 13398 14976 13404
rect 14936 12986 14964 13398
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 15120 12646 15148 14826
rect 15212 14346 15240 16050
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15212 12434 15240 13874
rect 15304 13841 15332 14758
rect 15396 14482 15424 14962
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15290 13832 15346 13841
rect 15290 13767 15346 13776
rect 15212 12406 15332 12434
rect 14922 12336 14978 12345
rect 14922 12271 14978 12280
rect 14936 11082 14964 12271
rect 15106 11792 15162 11801
rect 15106 11727 15162 11736
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 15120 8362 15148 11727
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14646 6896 14702 6905
rect 14646 6831 14702 6840
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14200 4282 14228 5306
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14200 4078 14228 4218
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14200 3058 14228 4014
rect 14568 3670 14596 4150
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14568 3126 14596 3606
rect 14660 3398 14688 6666
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14844 2922 14872 8230
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14924 5840 14976 5846
rect 14924 5782 14976 5788
rect 14936 3126 14964 5782
rect 15028 5370 15056 7414
rect 15212 6390 15240 10474
rect 15304 8090 15332 12406
rect 15396 10554 15424 14418
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 10849 15516 13670
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15580 11762 15608 13262
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15474 10840 15530 10849
rect 15474 10775 15530 10784
rect 15396 10526 15516 10554
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15396 9761 15424 10406
rect 15382 9752 15438 9761
rect 15382 9687 15438 9696
rect 15488 9382 15516 10526
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 10266 15608 10474
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15672 9654 15700 14282
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15382 6760 15438 6769
rect 15382 6695 15438 6704
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 15120 3602 15148 6054
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15212 4622 15240 5034
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15212 3602 15240 4558
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 15304 3058 15332 3878
rect 15396 3194 15424 6695
rect 15764 4554 15792 15846
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 13394 15884 14214
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 11286 15884 12038
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15842 10840 15898 10849
rect 15842 10775 15898 10784
rect 15856 10266 15884 10775
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15948 10146 15976 17138
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16316 15094 16344 16730
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16394 16008 16450 16017
rect 16394 15943 16450 15952
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 15856 10118 15976 10146
rect 15856 9926 15884 10118
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15856 8906 15884 9318
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15856 6798 15884 8842
rect 15948 8566 15976 9998
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 16040 6254 16068 14418
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 16132 10062 16160 13806
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16316 13161 16344 13194
rect 16302 13152 16358 13161
rect 16302 13087 16358 13096
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16224 10810 16252 12718
rect 16316 12374 16344 12922
rect 16408 12714 16436 15943
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16224 10470 16252 10746
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16408 9994 16436 10950
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15672 3466 15700 3946
rect 15750 3496 15806 3505
rect 15660 3460 15712 3466
rect 15750 3431 15752 3440
rect 15660 3402 15712 3408
rect 15804 3431 15806 3440
rect 15752 3402 15804 3408
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 13912 2848 13964 2854
rect 16132 2836 16160 9658
rect 16224 2990 16252 9862
rect 16408 9722 16436 9930
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16316 2990 16344 7958
rect 16394 7440 16450 7449
rect 16394 7375 16450 7384
rect 16408 6866 16436 7375
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16500 3194 16528 16390
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16592 16017 16620 16050
rect 16578 16008 16634 16017
rect 16578 15943 16634 15952
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16592 12782 16620 15846
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16592 7206 16620 12378
rect 16684 10742 16712 17138
rect 16950 16892 17258 16901
rect 16950 16890 16956 16892
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17252 16890 17258 16892
rect 17012 16838 17014 16890
rect 17194 16838 17196 16890
rect 16950 16836 16956 16838
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 17252 16836 17258 16838
rect 16950 16827 17258 16836
rect 18064 16794 18092 19200
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16776 14906 16804 16118
rect 16868 15706 16896 16458
rect 16950 15804 17258 15813
rect 16950 15802 16956 15804
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17252 15802 17258 15804
rect 17012 15750 17014 15802
rect 17194 15750 17196 15802
rect 16950 15748 16956 15750
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 17252 15748 17258 15750
rect 16950 15739 17258 15748
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16946 14920 17002 14929
rect 16776 14878 16896 14906
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16776 13433 16804 14758
rect 16762 13424 16818 13433
rect 16762 13359 16818 13368
rect 16868 12753 16896 14878
rect 16946 14855 16948 14864
rect 17000 14855 17002 14864
rect 16948 14826 17000 14832
rect 16950 14716 17258 14725
rect 16950 14714 16956 14716
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17252 14714 17258 14716
rect 17012 14662 17014 14714
rect 17194 14662 17196 14714
rect 16950 14660 16956 14662
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 17252 14660 17258 14662
rect 16950 14651 17258 14660
rect 16950 13628 17258 13637
rect 16950 13626 16956 13628
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17252 13626 17258 13628
rect 17012 13574 17014 13626
rect 17194 13574 17196 13626
rect 16950 13572 16956 13574
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 17252 13572 17258 13574
rect 16950 13563 17258 13572
rect 16854 12744 16910 12753
rect 16854 12679 16910 12688
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16776 12442 16804 12582
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16762 12336 16818 12345
rect 16762 12271 16818 12280
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16684 5386 16712 10542
rect 16776 6730 16804 12271
rect 16868 11218 16896 12582
rect 16950 12540 17258 12549
rect 16950 12538 16956 12540
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17252 12538 17258 12540
rect 17012 12486 17014 12538
rect 17194 12486 17196 12538
rect 16950 12484 16956 12486
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 17252 12484 17258 12486
rect 16950 12475 17258 12484
rect 17328 12434 17356 16526
rect 17610 16348 17918 16357
rect 17610 16346 17616 16348
rect 17672 16346 17696 16348
rect 17752 16346 17776 16348
rect 17832 16346 17856 16348
rect 17912 16346 17918 16348
rect 17672 16294 17674 16346
rect 17854 16294 17856 16346
rect 17610 16292 17616 16294
rect 17672 16292 17696 16294
rect 17752 16292 17776 16294
rect 17832 16292 17856 16294
rect 17912 16292 17918 16294
rect 17610 16283 17918 16292
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17236 12406 17356 12434
rect 17236 11558 17264 12406
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 16950 11452 17258 11461
rect 16950 11450 16956 11452
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17252 11450 17258 11452
rect 17012 11398 17014 11450
rect 17194 11398 17196 11450
rect 16950 11396 16956 11398
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 17252 11396 17258 11398
rect 16950 11387 17258 11396
rect 17130 11248 17186 11257
rect 16856 11212 16908 11218
rect 17130 11183 17186 11192
rect 16856 11154 16908 11160
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 16868 10198 16896 10678
rect 16960 10606 16988 11086
rect 17144 10810 17172 11183
rect 17328 11098 17356 12310
rect 17236 11070 17356 11098
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17236 10742 17264 11070
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17236 10606 17264 10678
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 16950 10364 17258 10373
rect 16950 10362 16956 10364
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17252 10362 17258 10364
rect 17012 10310 17014 10362
rect 17194 10310 17196 10362
rect 16950 10308 16956 10310
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 17252 10308 17258 10310
rect 16950 10299 17258 10308
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16960 9674 16988 10066
rect 16868 9646 16988 9674
rect 16868 7342 16896 9646
rect 16950 9276 17258 9285
rect 16950 9274 16956 9276
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17252 9274 17258 9276
rect 17012 9222 17014 9274
rect 17194 9222 17196 9274
rect 16950 9220 16956 9222
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 17252 9220 17258 9222
rect 16950 9211 17258 9220
rect 16950 8188 17258 8197
rect 16950 8186 16956 8188
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17252 8186 17258 8188
rect 17012 8134 17014 8186
rect 17194 8134 17196 8186
rect 16950 8132 16956 8134
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 17252 8132 17258 8134
rect 16950 8123 17258 8132
rect 17328 7818 17356 10950
rect 17420 9625 17448 15846
rect 17512 11014 17540 15982
rect 17610 15260 17918 15269
rect 17610 15258 17616 15260
rect 17672 15258 17696 15260
rect 17752 15258 17776 15260
rect 17832 15258 17856 15260
rect 17912 15258 17918 15260
rect 17672 15206 17674 15258
rect 17854 15206 17856 15258
rect 17610 15204 17616 15206
rect 17672 15204 17696 15206
rect 17752 15204 17776 15206
rect 17832 15204 17856 15206
rect 17912 15204 17918 15206
rect 17610 15195 17918 15204
rect 17610 14172 17918 14181
rect 17610 14170 17616 14172
rect 17672 14170 17696 14172
rect 17752 14170 17776 14172
rect 17832 14170 17856 14172
rect 17912 14170 17918 14172
rect 17672 14118 17674 14170
rect 17854 14118 17856 14170
rect 17610 14116 17616 14118
rect 17672 14116 17696 14118
rect 17752 14116 17776 14118
rect 17832 14116 17856 14118
rect 17912 14116 17918 14118
rect 17610 14107 17918 14116
rect 17610 13084 17918 13093
rect 17610 13082 17616 13084
rect 17672 13082 17696 13084
rect 17752 13082 17776 13084
rect 17832 13082 17856 13084
rect 17912 13082 17918 13084
rect 17672 13030 17674 13082
rect 17854 13030 17856 13082
rect 17610 13028 17616 13030
rect 17672 13028 17696 13030
rect 17752 13028 17776 13030
rect 17832 13028 17856 13030
rect 17912 13028 17918 13030
rect 17610 13019 17918 13028
rect 17610 11996 17918 12005
rect 17610 11994 17616 11996
rect 17672 11994 17696 11996
rect 17752 11994 17776 11996
rect 17832 11994 17856 11996
rect 17912 11994 17918 11996
rect 17672 11942 17674 11994
rect 17854 11942 17856 11994
rect 17610 11940 17616 11942
rect 17672 11940 17696 11942
rect 17752 11940 17776 11942
rect 17832 11940 17856 11942
rect 17912 11940 17918 11942
rect 17610 11931 17918 11940
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17610 10908 17918 10917
rect 17610 10906 17616 10908
rect 17672 10906 17696 10908
rect 17752 10906 17776 10908
rect 17832 10906 17856 10908
rect 17912 10906 17918 10908
rect 17672 10854 17674 10906
rect 17854 10854 17856 10906
rect 17610 10852 17616 10854
rect 17672 10852 17696 10854
rect 17752 10852 17776 10854
rect 17832 10852 17856 10854
rect 17912 10852 17918 10854
rect 17610 10843 17918 10852
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17512 10538 17540 10678
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17500 10532 17552 10538
rect 17500 10474 17552 10480
rect 17406 9616 17462 9625
rect 17406 9551 17462 9560
rect 17316 7812 17368 7818
rect 17316 7754 17368 7760
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16868 5574 16896 7278
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 16950 7100 17258 7109
rect 16950 7098 16956 7100
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17252 7098 17258 7100
rect 17012 7046 17014 7098
rect 17194 7046 17196 7098
rect 16950 7044 16956 7046
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 17252 7044 17258 7046
rect 16950 7035 17258 7044
rect 16950 6012 17258 6021
rect 16950 6010 16956 6012
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17252 6010 17258 6012
rect 17012 5958 17014 6010
rect 17194 5958 17196 6010
rect 16950 5956 16956 5958
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 17252 5956 17258 5958
rect 16950 5947 17258 5956
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16684 5358 16896 5386
rect 16762 5264 16818 5273
rect 16762 5199 16818 5208
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16776 3058 16804 5199
rect 16868 4826 16896 5358
rect 16950 4924 17258 4933
rect 16950 4922 16956 4924
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17252 4922 17258 4924
rect 17012 4870 17014 4922
rect 17194 4870 17196 4922
rect 16950 4868 16956 4870
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 17252 4868 17258 4870
rect 16950 4859 17258 4868
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16950 3836 17258 3845
rect 16950 3834 16956 3836
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17252 3834 17258 3836
rect 17012 3782 17014 3834
rect 17194 3782 17196 3834
rect 16950 3780 16956 3782
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 17252 3780 17258 3782
rect 16950 3771 17258 3780
rect 17328 3466 17356 7142
rect 17420 5030 17448 7346
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17316 3460 17368 3466
rect 17316 3402 17368 3408
rect 17420 3058 17448 4762
rect 17512 4282 17540 10474
rect 17604 10130 17632 10542
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17696 10062 17724 10746
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17610 9820 17918 9829
rect 17610 9818 17616 9820
rect 17672 9818 17696 9820
rect 17752 9818 17776 9820
rect 17832 9818 17856 9820
rect 17912 9818 17918 9820
rect 17672 9766 17674 9818
rect 17854 9766 17856 9818
rect 17610 9764 17616 9766
rect 17672 9764 17696 9766
rect 17752 9764 17776 9766
rect 17832 9764 17856 9766
rect 17912 9764 17918 9766
rect 17610 9755 17918 9764
rect 17610 8732 17918 8741
rect 17610 8730 17616 8732
rect 17672 8730 17696 8732
rect 17752 8730 17776 8732
rect 17832 8730 17856 8732
rect 17912 8730 17918 8732
rect 17672 8678 17674 8730
rect 17854 8678 17856 8730
rect 17610 8676 17616 8678
rect 17672 8676 17696 8678
rect 17752 8676 17776 8678
rect 17832 8676 17856 8678
rect 17912 8676 17918 8678
rect 17610 8667 17918 8676
rect 17610 7644 17918 7653
rect 17610 7642 17616 7644
rect 17672 7642 17696 7644
rect 17752 7642 17776 7644
rect 17832 7642 17856 7644
rect 17912 7642 17918 7644
rect 17672 7590 17674 7642
rect 17854 7590 17856 7642
rect 17610 7588 17616 7590
rect 17672 7588 17696 7590
rect 17752 7588 17776 7590
rect 17832 7588 17856 7590
rect 17912 7588 17918 7590
rect 17610 7579 17918 7588
rect 17610 6556 17918 6565
rect 17610 6554 17616 6556
rect 17672 6554 17696 6556
rect 17752 6554 17776 6556
rect 17832 6554 17856 6556
rect 17912 6554 17918 6556
rect 17672 6502 17674 6554
rect 17854 6502 17856 6554
rect 17610 6500 17616 6502
rect 17672 6500 17696 6502
rect 17752 6500 17776 6502
rect 17832 6500 17856 6502
rect 17912 6500 17918 6502
rect 17610 6491 17918 6500
rect 17972 6361 18000 16662
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 18064 11642 18092 15846
rect 18156 12986 18184 15914
rect 18248 15745 18276 16050
rect 18234 15736 18290 15745
rect 18234 15671 18290 15680
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18156 12345 18184 12786
rect 18432 12434 18460 12922
rect 18432 12406 18644 12434
rect 18142 12336 18198 12345
rect 18142 12271 18198 12280
rect 18064 11614 18460 11642
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18156 10470 18184 11494
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17958 6352 18014 6361
rect 18064 6322 18092 9998
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 18156 9625 18184 9930
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18142 9616 18198 9625
rect 18142 9551 18198 9560
rect 18248 8974 18276 9862
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 17958 6287 18014 6296
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 18156 5710 18184 8298
rect 18340 7857 18368 10406
rect 18432 9674 18460 11614
rect 18432 9646 18552 9674
rect 18326 7848 18382 7857
rect 18326 7783 18382 7792
rect 18418 6216 18474 6225
rect 18418 6151 18420 6160
rect 18472 6151 18474 6160
rect 18420 6122 18472 6128
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17610 5468 17918 5477
rect 17610 5466 17616 5468
rect 17672 5466 17696 5468
rect 17752 5466 17776 5468
rect 17832 5466 17856 5468
rect 17912 5466 17918 5468
rect 17672 5414 17674 5466
rect 17854 5414 17856 5466
rect 17610 5412 17616 5414
rect 17672 5412 17696 5414
rect 17752 5412 17776 5414
rect 17832 5412 17856 5414
rect 17912 5412 17918 5414
rect 17610 5403 17918 5412
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17880 4570 17908 4966
rect 17880 4542 18000 4570
rect 17610 4380 17918 4389
rect 17610 4378 17616 4380
rect 17672 4378 17696 4380
rect 17752 4378 17776 4380
rect 17832 4378 17856 4380
rect 17912 4378 17918 4380
rect 17672 4326 17674 4378
rect 17854 4326 17856 4378
rect 17610 4324 17616 4326
rect 17672 4324 17696 4326
rect 17752 4324 17776 4326
rect 17832 4324 17856 4326
rect 17912 4324 17918 4326
rect 17610 4315 17918 4324
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17972 4162 18000 4542
rect 18064 4214 18092 5510
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 17880 4134 18000 4162
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 17592 4072 17644 4078
rect 17498 4040 17554 4049
rect 17592 4014 17644 4020
rect 17498 3975 17554 3984
rect 17512 3738 17540 3975
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17604 3618 17632 4014
rect 17512 3590 17632 3618
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 17512 2922 17540 3590
rect 17880 3534 17908 4134
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18156 3738 18184 3946
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18142 3496 18198 3505
rect 18142 3431 18144 3440
rect 18196 3431 18198 3440
rect 18144 3402 18196 3408
rect 17610 3292 17918 3301
rect 17610 3290 17616 3292
rect 17672 3290 17696 3292
rect 17752 3290 17776 3292
rect 17832 3290 17856 3292
rect 17912 3290 17918 3292
rect 17672 3238 17674 3290
rect 17854 3238 17856 3290
rect 17610 3236 17616 3238
rect 17672 3236 17696 3238
rect 17752 3236 17776 3238
rect 17832 3236 17856 3238
rect 17912 3236 17918 3238
rect 17610 3227 17918 3236
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 16304 2848 16356 2854
rect 16132 2808 16304 2836
rect 13912 2790 13964 2796
rect 16304 2790 16356 2796
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 16316 2582 16344 2790
rect 16950 2748 17258 2757
rect 16950 2746 16956 2748
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17252 2746 17258 2748
rect 17012 2694 17014 2746
rect 17194 2694 17196 2746
rect 16950 2692 16956 2694
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 17252 2692 17258 2694
rect 16950 2683 17258 2692
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 17604 2446 17632 3062
rect 18340 2650 18368 5238
rect 18432 4282 18460 5578
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18524 3602 18552 9646
rect 18616 3942 18644 12406
rect 18708 10742 18736 14894
rect 18696 10736 18748 10742
rect 18696 10678 18748 10684
rect 18708 4078 18736 10678
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18616 3670 18644 3878
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18800 2990 18828 10474
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 14200 800 14228 2246
rect 17420 800 17448 2246
rect 17610 2204 17918 2213
rect 17610 2202 17616 2204
rect 17672 2202 17696 2204
rect 17752 2202 17776 2204
rect 17832 2202 17856 2204
rect 17912 2202 17918 2204
rect 17672 2150 17674 2202
rect 17854 2150 17856 2202
rect 17610 2148 17616 2150
rect 17672 2148 17696 2150
rect 17752 2148 17776 2150
rect 17832 2148 17856 2150
rect 17912 2148 17918 2150
rect 17610 2139 17918 2148
rect 17972 1986 18000 2382
rect 17880 1958 18000 1986
rect 18 0 74 800
rect 2594 0 2650 800
rect 5814 0 5870 800
rect 8390 0 8446 800
rect 11610 0 11666 800
rect 14186 0 14242 800
rect 17406 0 17462 800
rect 17880 105 17908 1958
rect 17866 96 17922 105
rect 17866 31 17922 40
<< via2 >>
rect 1582 18400 1638 18456
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 7616 17434 7672 17436
rect 7696 17434 7752 17436
rect 7776 17434 7832 17436
rect 7856 17434 7912 17436
rect 7616 17382 7662 17434
rect 7662 17382 7672 17434
rect 7696 17382 7726 17434
rect 7726 17382 7738 17434
rect 7738 17382 7752 17434
rect 7776 17382 7790 17434
rect 7790 17382 7802 17434
rect 7802 17382 7832 17434
rect 7856 17382 7866 17434
rect 7866 17382 7912 17434
rect 7616 17380 7672 17382
rect 7696 17380 7752 17382
rect 7776 17380 7832 17382
rect 7856 17380 7912 17382
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 1490 15952 1546 16008
rect 3238 16088 3294 16144
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 1582 15000 1638 15056
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 2502 13932 2558 13968
rect 2502 13912 2504 13932
rect 2504 13912 2556 13932
rect 2556 13912 2558 13932
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 2134 12824 2190 12880
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 1582 12280 1638 12336
rect 1950 11756 2006 11792
rect 1950 11736 1952 11756
rect 1952 11736 2004 11756
rect 2004 11736 2006 11756
rect 2226 11736 2282 11792
rect 1766 11192 1822 11248
rect 938 8880 994 8936
rect 938 6160 994 6216
rect 1582 5616 1638 5672
rect 1398 3440 1454 3496
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1950 6160 2006 6216
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2042 5108 2044 5128
rect 2044 5108 2096 5128
rect 2096 5108 2098 5128
rect 2042 5072 2098 5108
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2134 4156 2136 4176
rect 2136 4156 2188 4176
rect 2188 4156 2190 4176
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 2870 12180 2872 12200
rect 2872 12180 2924 12200
rect 2924 12180 2926 12200
rect 2870 12144 2926 12180
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 3054 12300 3110 12336
rect 3054 12280 3056 12300
rect 3056 12280 3108 12300
rect 3108 12280 3110 12300
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 2502 10512 2558 10568
rect 2502 10240 2558 10296
rect 2410 5208 2466 5264
rect 2134 4120 2190 4156
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3054 9968 3110 10024
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 3422 14320 3478 14376
rect 3054 5480 3110 5536
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 4066 16088 4122 16144
rect 3974 15544 4030 15600
rect 3882 11092 3884 11112
rect 3884 11092 3936 11112
rect 3936 11092 3938 11112
rect 3882 11056 3938 11092
rect 3698 7928 3754 7984
rect 3698 7248 3754 7304
rect 3606 5480 3662 5536
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 3790 6840 3846 6896
rect 4066 13776 4122 13832
rect 5354 16632 5410 16688
rect 4342 13812 4344 13832
rect 4344 13812 4396 13832
rect 4396 13812 4398 13832
rect 4342 13776 4398 13812
rect 5170 15308 5172 15328
rect 5172 15308 5224 15328
rect 5224 15308 5226 15328
rect 5170 15272 5226 15308
rect 4802 14456 4858 14512
rect 4158 12144 4214 12200
rect 4526 12688 4582 12744
rect 4434 10648 4490 10704
rect 4250 5480 4306 5536
rect 4250 4664 4306 4720
rect 4342 3984 4398 4040
rect 5170 13368 5226 13424
rect 5078 10920 5134 10976
rect 5354 12144 5410 12200
rect 5262 10240 5318 10296
rect 5170 9580 5226 9616
rect 5170 9560 5172 9580
rect 5172 9560 5224 9580
rect 5224 9560 5226 9580
rect 4986 5072 5042 5128
rect 5538 9016 5594 9072
rect 5262 4820 5318 4856
rect 5262 4800 5264 4820
rect 5264 4800 5316 4820
rect 5316 4800 5318 4820
rect 5722 8472 5778 8528
rect 6090 11736 6146 11792
rect 5722 7112 5778 7168
rect 5722 6840 5778 6896
rect 5630 6024 5686 6080
rect 5814 6740 5816 6760
rect 5816 6740 5868 6760
rect 5868 6740 5870 6760
rect 5814 6704 5870 6740
rect 6090 9424 6146 9480
rect 5998 7656 6054 7712
rect 6366 13912 6422 13968
rect 6366 12824 6422 12880
rect 6956 16890 7012 16892
rect 7036 16890 7092 16892
rect 7116 16890 7172 16892
rect 7196 16890 7252 16892
rect 6956 16838 7002 16890
rect 7002 16838 7012 16890
rect 7036 16838 7066 16890
rect 7066 16838 7078 16890
rect 7078 16838 7092 16890
rect 7116 16838 7130 16890
rect 7130 16838 7142 16890
rect 7142 16838 7172 16890
rect 7196 16838 7206 16890
rect 7206 16838 7252 16890
rect 6956 16836 7012 16838
rect 7036 16836 7092 16838
rect 7116 16836 7172 16838
rect 7196 16836 7252 16838
rect 7616 16346 7672 16348
rect 7696 16346 7752 16348
rect 7776 16346 7832 16348
rect 7856 16346 7912 16348
rect 7616 16294 7662 16346
rect 7662 16294 7672 16346
rect 7696 16294 7726 16346
rect 7726 16294 7738 16346
rect 7738 16294 7752 16346
rect 7776 16294 7790 16346
rect 7790 16294 7802 16346
rect 7802 16294 7832 16346
rect 7856 16294 7866 16346
rect 7866 16294 7912 16346
rect 7616 16292 7672 16294
rect 7696 16292 7752 16294
rect 7776 16292 7832 16294
rect 7856 16292 7912 16294
rect 6734 15408 6790 15464
rect 6550 11636 6552 11656
rect 6552 11636 6604 11656
rect 6604 11636 6606 11656
rect 6550 11600 6606 11636
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 7378 15952 7434 16008
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 6274 7520 6330 7576
rect 6090 5480 6146 5536
rect 4342 3032 4398 3088
rect 5170 3032 5226 3088
rect 938 2796 940 2816
rect 940 2796 992 2816
rect 992 2796 994 2816
rect 938 2760 994 2796
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 6090 4528 6146 4584
rect 6550 7656 6606 7712
rect 6734 7656 6790 7712
rect 6550 6976 6606 7032
rect 6734 7112 6790 7168
rect 6734 6840 6790 6896
rect 6642 6296 6698 6352
rect 6642 6024 6698 6080
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 6918 9424 6974 9480
rect 7194 9696 7250 9752
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 7746 12416 7802 12472
rect 8666 15000 8722 15056
rect 8206 13776 8262 13832
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 7654 11620 7710 11656
rect 7654 11600 7656 11620
rect 7656 11600 7708 11620
rect 7708 11600 7710 11620
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 8114 11600 8170 11656
rect 8482 12280 8538 12336
rect 8482 10648 8538 10704
rect 8298 9832 8354 9888
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 7470 9288 7526 9344
rect 7470 9152 7526 9208
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 6918 7520 6974 7576
rect 7102 7792 7158 7848
rect 7286 7792 7342 7848
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 6826 5752 6882 5808
rect 9126 15272 9182 15328
rect 8574 9968 8630 10024
rect 8850 11056 8906 11112
rect 8666 9696 8722 9752
rect 7930 9560 7986 9616
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 8206 8608 8262 8664
rect 8206 7248 8262 7304
rect 8390 7928 8446 7984
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 7838 5888 7894 5944
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 7654 5244 7656 5264
rect 7656 5244 7708 5264
rect 7708 5244 7710 5264
rect 7654 5208 7710 5244
rect 7654 4820 7710 4856
rect 7654 4800 7656 4820
rect 7656 4800 7708 4820
rect 7708 4800 7710 4820
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 6550 2896 6606 2952
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 8298 6160 8354 6216
rect 8206 4664 8262 4720
rect 8758 6568 8814 6624
rect 8758 6024 8814 6080
rect 8666 5888 8722 5944
rect 8298 2896 8354 2952
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 9126 11056 9182 11112
rect 9402 8472 9458 8528
rect 9402 5072 9458 5128
rect 9310 4120 9366 4176
rect 9126 2524 9128 2544
rect 9128 2524 9180 2544
rect 9180 2524 9182 2544
rect 9126 2488 9182 2524
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 9770 11464 9826 11520
rect 9678 11328 9734 11384
rect 10046 11872 10102 11928
rect 9862 8064 9918 8120
rect 9678 4684 9734 4720
rect 9678 4664 9680 4684
rect 9680 4664 9732 4684
rect 9732 4664 9734 4684
rect 9586 3576 9642 3632
rect 10322 14184 10378 14240
rect 10230 12280 10286 12336
rect 10598 15272 10654 15328
rect 10782 15136 10838 15192
rect 10690 14728 10746 14784
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 17866 18400 17922 18456
rect 17616 17434 17672 17436
rect 17696 17434 17752 17436
rect 17776 17434 17832 17436
rect 17856 17434 17912 17436
rect 17616 17382 17662 17434
rect 17662 17382 17672 17434
rect 17696 17382 17726 17434
rect 17726 17382 17738 17434
rect 17738 17382 17752 17434
rect 17776 17382 17790 17434
rect 17790 17382 17802 17434
rect 17802 17382 17832 17434
rect 17856 17382 17866 17434
rect 17866 17382 17912 17434
rect 17616 17380 17672 17382
rect 17696 17380 17752 17382
rect 17776 17380 17832 17382
rect 17856 17380 17912 17382
rect 11956 16890 12012 16892
rect 12036 16890 12092 16892
rect 12116 16890 12172 16892
rect 12196 16890 12252 16892
rect 11956 16838 12002 16890
rect 12002 16838 12012 16890
rect 12036 16838 12066 16890
rect 12066 16838 12078 16890
rect 12078 16838 12092 16890
rect 12116 16838 12130 16890
rect 12130 16838 12142 16890
rect 12142 16838 12172 16890
rect 12196 16838 12206 16890
rect 12206 16838 12252 16890
rect 11956 16836 12012 16838
rect 12036 16836 12092 16838
rect 12116 16836 12172 16838
rect 12196 16836 12252 16838
rect 10414 11328 10470 11384
rect 10230 11056 10286 11112
rect 10230 10920 10286 10976
rect 10598 11464 10654 11520
rect 10506 9424 10562 9480
rect 9954 4564 9956 4584
rect 9956 4564 10008 4584
rect 10008 4564 10010 4584
rect 9954 4528 10010 4564
rect 10138 4528 10194 4584
rect 11150 15544 11206 15600
rect 13174 16496 13230 16552
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 12622 16088 12678 16144
rect 12806 16088 12862 16144
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 11978 15544 12034 15600
rect 11426 14356 11428 14376
rect 11428 14356 11480 14376
rect 11480 14356 11482 14376
rect 11426 14320 11482 14356
rect 11610 14728 11666 14784
rect 11886 15156 11942 15192
rect 11886 15136 11888 15156
rect 11888 15136 11940 15156
rect 11940 15136 11942 15156
rect 12438 15272 12494 15328
rect 12162 15000 12218 15056
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 11978 14476 12034 14512
rect 11978 14456 11980 14476
rect 11980 14456 12032 14476
rect 12032 14456 12034 14476
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 11058 11348 11114 11384
rect 11058 11328 11060 11348
rect 11060 11328 11112 11348
rect 11112 11328 11114 11348
rect 11058 11192 11114 11248
rect 10966 11056 11022 11112
rect 11242 10104 11298 10160
rect 10874 5072 10930 5128
rect 11058 6704 11114 6760
rect 10782 3984 10838 4040
rect 11150 3712 11206 3768
rect 12254 12824 12310 12880
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 11886 11872 11942 11928
rect 11426 6432 11482 6488
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 12254 11228 12256 11248
rect 12256 11228 12308 11248
rect 12308 11228 12310 11248
rect 12254 11192 12310 11228
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 12622 15816 12678 15872
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 13266 15816 13322 15872
rect 12898 14320 12954 14376
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 12990 12688 13046 12744
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 12530 10104 12586 10160
rect 12438 9424 12494 9480
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 11702 6704 11758 6760
rect 11610 6432 11666 6488
rect 11426 4800 11482 4856
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 11886 4684 11942 4720
rect 11886 4664 11888 4684
rect 11888 4664 11940 4684
rect 11940 4664 11942 4684
rect 11794 3848 11850 3904
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 11886 3476 11888 3496
rect 11888 3476 11940 3496
rect 11940 3476 11942 3496
rect 11886 3440 11942 3476
rect 12162 3168 12218 3224
rect 12346 3168 12402 3224
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 12070 3032 12126 3088
rect 11794 2896 11850 2952
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 12530 3032 12586 3088
rect 13358 11600 13414 11656
rect 13358 10648 13414 10704
rect 13910 15272 13966 15328
rect 13818 13252 13874 13288
rect 13818 13232 13820 13252
rect 13820 13232 13872 13252
rect 13872 13232 13874 13252
rect 14830 16088 14886 16144
rect 14278 15544 14334 15600
rect 14370 15428 14426 15464
rect 14370 15408 14372 15428
rect 14372 15408 14424 15428
rect 14424 15408 14426 15428
rect 13634 10512 13690 10568
rect 13450 8472 13506 8528
rect 13634 10240 13690 10296
rect 13542 8200 13598 8256
rect 14094 12180 14096 12200
rect 14096 12180 14148 12200
rect 14148 12180 14150 12200
rect 14094 12144 14150 12180
rect 13818 8472 13874 8528
rect 13818 6160 13874 6216
rect 13726 5072 13782 5128
rect 15014 15272 15070 15328
rect 15290 13776 15346 13832
rect 14922 12280 14978 12336
rect 15106 11736 15162 11792
rect 14646 6840 14702 6896
rect 15474 10784 15530 10840
rect 15382 9696 15438 9752
rect 15382 6704 15438 6760
rect 15842 10784 15898 10840
rect 16394 15952 16450 16008
rect 16302 13096 16358 13152
rect 15750 3460 15806 3496
rect 15750 3440 15752 3460
rect 15752 3440 15804 3460
rect 15804 3440 15806 3460
rect 16394 7384 16450 7440
rect 16578 15952 16634 16008
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 17002 16890
rect 17002 16838 17012 16890
rect 17036 16838 17066 16890
rect 17066 16838 17078 16890
rect 17078 16838 17092 16890
rect 17116 16838 17130 16890
rect 17130 16838 17142 16890
rect 17142 16838 17172 16890
rect 17196 16838 17206 16890
rect 17206 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 17002 15802
rect 17002 15750 17012 15802
rect 17036 15750 17066 15802
rect 17066 15750 17078 15802
rect 17078 15750 17092 15802
rect 17116 15750 17130 15802
rect 17130 15750 17142 15802
rect 17142 15750 17172 15802
rect 17196 15750 17206 15802
rect 17206 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16762 13368 16818 13424
rect 16946 14884 17002 14920
rect 16946 14864 16948 14884
rect 16948 14864 17000 14884
rect 17000 14864 17002 14884
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 17002 14714
rect 17002 14662 17012 14714
rect 17036 14662 17066 14714
rect 17066 14662 17078 14714
rect 17078 14662 17092 14714
rect 17116 14662 17130 14714
rect 17130 14662 17142 14714
rect 17142 14662 17172 14714
rect 17196 14662 17206 14714
rect 17206 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 17002 13626
rect 17002 13574 17012 13626
rect 17036 13574 17066 13626
rect 17066 13574 17078 13626
rect 17078 13574 17092 13626
rect 17116 13574 17130 13626
rect 17130 13574 17142 13626
rect 17142 13574 17172 13626
rect 17196 13574 17206 13626
rect 17206 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16854 12688 16910 12744
rect 16762 12280 16818 12336
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 17002 12538
rect 17002 12486 17012 12538
rect 17036 12486 17066 12538
rect 17066 12486 17078 12538
rect 17078 12486 17092 12538
rect 17116 12486 17130 12538
rect 17130 12486 17142 12538
rect 17142 12486 17172 12538
rect 17196 12486 17206 12538
rect 17206 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 17616 16346 17672 16348
rect 17696 16346 17752 16348
rect 17776 16346 17832 16348
rect 17856 16346 17912 16348
rect 17616 16294 17662 16346
rect 17662 16294 17672 16346
rect 17696 16294 17726 16346
rect 17726 16294 17738 16346
rect 17738 16294 17752 16346
rect 17776 16294 17790 16346
rect 17790 16294 17802 16346
rect 17802 16294 17832 16346
rect 17856 16294 17866 16346
rect 17866 16294 17912 16346
rect 17616 16292 17672 16294
rect 17696 16292 17752 16294
rect 17776 16292 17832 16294
rect 17856 16292 17912 16294
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 17002 11450
rect 17002 11398 17012 11450
rect 17036 11398 17066 11450
rect 17066 11398 17078 11450
rect 17078 11398 17092 11450
rect 17116 11398 17130 11450
rect 17130 11398 17142 11450
rect 17142 11398 17172 11450
rect 17196 11398 17206 11450
rect 17206 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 17130 11192 17186 11248
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 17002 10362
rect 17002 10310 17012 10362
rect 17036 10310 17066 10362
rect 17066 10310 17078 10362
rect 17078 10310 17092 10362
rect 17116 10310 17130 10362
rect 17130 10310 17142 10362
rect 17142 10310 17172 10362
rect 17196 10310 17206 10362
rect 17206 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 17002 9274
rect 17002 9222 17012 9274
rect 17036 9222 17066 9274
rect 17066 9222 17078 9274
rect 17078 9222 17092 9274
rect 17116 9222 17130 9274
rect 17130 9222 17142 9274
rect 17142 9222 17172 9274
rect 17196 9222 17206 9274
rect 17206 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 17002 8186
rect 17002 8134 17012 8186
rect 17036 8134 17066 8186
rect 17066 8134 17078 8186
rect 17078 8134 17092 8186
rect 17116 8134 17130 8186
rect 17130 8134 17142 8186
rect 17142 8134 17172 8186
rect 17196 8134 17206 8186
rect 17206 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 17616 15258 17672 15260
rect 17696 15258 17752 15260
rect 17776 15258 17832 15260
rect 17856 15258 17912 15260
rect 17616 15206 17662 15258
rect 17662 15206 17672 15258
rect 17696 15206 17726 15258
rect 17726 15206 17738 15258
rect 17738 15206 17752 15258
rect 17776 15206 17790 15258
rect 17790 15206 17802 15258
rect 17802 15206 17832 15258
rect 17856 15206 17866 15258
rect 17866 15206 17912 15258
rect 17616 15204 17672 15206
rect 17696 15204 17752 15206
rect 17776 15204 17832 15206
rect 17856 15204 17912 15206
rect 17616 14170 17672 14172
rect 17696 14170 17752 14172
rect 17776 14170 17832 14172
rect 17856 14170 17912 14172
rect 17616 14118 17662 14170
rect 17662 14118 17672 14170
rect 17696 14118 17726 14170
rect 17726 14118 17738 14170
rect 17738 14118 17752 14170
rect 17776 14118 17790 14170
rect 17790 14118 17802 14170
rect 17802 14118 17832 14170
rect 17856 14118 17866 14170
rect 17866 14118 17912 14170
rect 17616 14116 17672 14118
rect 17696 14116 17752 14118
rect 17776 14116 17832 14118
rect 17856 14116 17912 14118
rect 17616 13082 17672 13084
rect 17696 13082 17752 13084
rect 17776 13082 17832 13084
rect 17856 13082 17912 13084
rect 17616 13030 17662 13082
rect 17662 13030 17672 13082
rect 17696 13030 17726 13082
rect 17726 13030 17738 13082
rect 17738 13030 17752 13082
rect 17776 13030 17790 13082
rect 17790 13030 17802 13082
rect 17802 13030 17832 13082
rect 17856 13030 17866 13082
rect 17866 13030 17912 13082
rect 17616 13028 17672 13030
rect 17696 13028 17752 13030
rect 17776 13028 17832 13030
rect 17856 13028 17912 13030
rect 17616 11994 17672 11996
rect 17696 11994 17752 11996
rect 17776 11994 17832 11996
rect 17856 11994 17912 11996
rect 17616 11942 17662 11994
rect 17662 11942 17672 11994
rect 17696 11942 17726 11994
rect 17726 11942 17738 11994
rect 17738 11942 17752 11994
rect 17776 11942 17790 11994
rect 17790 11942 17802 11994
rect 17802 11942 17832 11994
rect 17856 11942 17866 11994
rect 17866 11942 17912 11994
rect 17616 11940 17672 11942
rect 17696 11940 17752 11942
rect 17776 11940 17832 11942
rect 17856 11940 17912 11942
rect 17616 10906 17672 10908
rect 17696 10906 17752 10908
rect 17776 10906 17832 10908
rect 17856 10906 17912 10908
rect 17616 10854 17662 10906
rect 17662 10854 17672 10906
rect 17696 10854 17726 10906
rect 17726 10854 17738 10906
rect 17738 10854 17752 10906
rect 17776 10854 17790 10906
rect 17790 10854 17802 10906
rect 17802 10854 17832 10906
rect 17856 10854 17866 10906
rect 17866 10854 17912 10906
rect 17616 10852 17672 10854
rect 17696 10852 17752 10854
rect 17776 10852 17832 10854
rect 17856 10852 17912 10854
rect 17406 9560 17462 9616
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 17002 7098
rect 17002 7046 17012 7098
rect 17036 7046 17066 7098
rect 17066 7046 17078 7098
rect 17078 7046 17092 7098
rect 17116 7046 17130 7098
rect 17130 7046 17142 7098
rect 17142 7046 17172 7098
rect 17196 7046 17206 7098
rect 17206 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 17002 6010
rect 17002 5958 17012 6010
rect 17036 5958 17066 6010
rect 17066 5958 17078 6010
rect 17078 5958 17092 6010
rect 17116 5958 17130 6010
rect 17130 5958 17142 6010
rect 17142 5958 17172 6010
rect 17196 5958 17206 6010
rect 17206 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16762 5208 16818 5264
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 17002 4922
rect 17002 4870 17012 4922
rect 17036 4870 17066 4922
rect 17066 4870 17078 4922
rect 17078 4870 17092 4922
rect 17116 4870 17130 4922
rect 17130 4870 17142 4922
rect 17142 4870 17172 4922
rect 17196 4870 17206 4922
rect 17206 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 17002 3834
rect 17002 3782 17012 3834
rect 17036 3782 17066 3834
rect 17066 3782 17078 3834
rect 17078 3782 17092 3834
rect 17116 3782 17130 3834
rect 17130 3782 17142 3834
rect 17142 3782 17172 3834
rect 17196 3782 17206 3834
rect 17206 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 17616 9818 17672 9820
rect 17696 9818 17752 9820
rect 17776 9818 17832 9820
rect 17856 9818 17912 9820
rect 17616 9766 17662 9818
rect 17662 9766 17672 9818
rect 17696 9766 17726 9818
rect 17726 9766 17738 9818
rect 17738 9766 17752 9818
rect 17776 9766 17790 9818
rect 17790 9766 17802 9818
rect 17802 9766 17832 9818
rect 17856 9766 17866 9818
rect 17866 9766 17912 9818
rect 17616 9764 17672 9766
rect 17696 9764 17752 9766
rect 17776 9764 17832 9766
rect 17856 9764 17912 9766
rect 17616 8730 17672 8732
rect 17696 8730 17752 8732
rect 17776 8730 17832 8732
rect 17856 8730 17912 8732
rect 17616 8678 17662 8730
rect 17662 8678 17672 8730
rect 17696 8678 17726 8730
rect 17726 8678 17738 8730
rect 17738 8678 17752 8730
rect 17776 8678 17790 8730
rect 17790 8678 17802 8730
rect 17802 8678 17832 8730
rect 17856 8678 17866 8730
rect 17866 8678 17912 8730
rect 17616 8676 17672 8678
rect 17696 8676 17752 8678
rect 17776 8676 17832 8678
rect 17856 8676 17912 8678
rect 17616 7642 17672 7644
rect 17696 7642 17752 7644
rect 17776 7642 17832 7644
rect 17856 7642 17912 7644
rect 17616 7590 17662 7642
rect 17662 7590 17672 7642
rect 17696 7590 17726 7642
rect 17726 7590 17738 7642
rect 17738 7590 17752 7642
rect 17776 7590 17790 7642
rect 17790 7590 17802 7642
rect 17802 7590 17832 7642
rect 17856 7590 17866 7642
rect 17866 7590 17912 7642
rect 17616 7588 17672 7590
rect 17696 7588 17752 7590
rect 17776 7588 17832 7590
rect 17856 7588 17912 7590
rect 17616 6554 17672 6556
rect 17696 6554 17752 6556
rect 17776 6554 17832 6556
rect 17856 6554 17912 6556
rect 17616 6502 17662 6554
rect 17662 6502 17672 6554
rect 17696 6502 17726 6554
rect 17726 6502 17738 6554
rect 17738 6502 17752 6554
rect 17776 6502 17790 6554
rect 17790 6502 17802 6554
rect 17802 6502 17832 6554
rect 17856 6502 17866 6554
rect 17866 6502 17912 6554
rect 17616 6500 17672 6502
rect 17696 6500 17752 6502
rect 17776 6500 17832 6502
rect 17856 6500 17912 6502
rect 18234 15680 18290 15736
rect 18142 12280 18198 12336
rect 17958 6296 18014 6352
rect 18142 9560 18198 9616
rect 18326 7792 18382 7848
rect 18418 6180 18474 6216
rect 18418 6160 18420 6180
rect 18420 6160 18472 6180
rect 18472 6160 18474 6180
rect 17616 5466 17672 5468
rect 17696 5466 17752 5468
rect 17776 5466 17832 5468
rect 17856 5466 17912 5468
rect 17616 5414 17662 5466
rect 17662 5414 17672 5466
rect 17696 5414 17726 5466
rect 17726 5414 17738 5466
rect 17738 5414 17752 5466
rect 17776 5414 17790 5466
rect 17790 5414 17802 5466
rect 17802 5414 17832 5466
rect 17856 5414 17866 5466
rect 17866 5414 17912 5466
rect 17616 5412 17672 5414
rect 17696 5412 17752 5414
rect 17776 5412 17832 5414
rect 17856 5412 17912 5414
rect 17616 4378 17672 4380
rect 17696 4378 17752 4380
rect 17776 4378 17832 4380
rect 17856 4378 17912 4380
rect 17616 4326 17662 4378
rect 17662 4326 17672 4378
rect 17696 4326 17726 4378
rect 17726 4326 17738 4378
rect 17738 4326 17752 4378
rect 17776 4326 17790 4378
rect 17790 4326 17802 4378
rect 17802 4326 17832 4378
rect 17856 4326 17866 4378
rect 17866 4326 17912 4378
rect 17616 4324 17672 4326
rect 17696 4324 17752 4326
rect 17776 4324 17832 4326
rect 17856 4324 17912 4326
rect 17498 3984 17554 4040
rect 18142 3460 18198 3496
rect 18142 3440 18144 3460
rect 18144 3440 18196 3460
rect 18196 3440 18198 3460
rect 17616 3290 17672 3292
rect 17696 3290 17752 3292
rect 17776 3290 17832 3292
rect 17856 3290 17912 3292
rect 17616 3238 17662 3290
rect 17662 3238 17672 3290
rect 17696 3238 17726 3290
rect 17726 3238 17738 3290
rect 17738 3238 17752 3290
rect 17776 3238 17790 3290
rect 17790 3238 17802 3290
rect 17802 3238 17832 3290
rect 17856 3238 17866 3290
rect 17866 3238 17912 3290
rect 17616 3236 17672 3238
rect 17696 3236 17752 3238
rect 17776 3236 17832 3238
rect 17856 3236 17912 3238
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 17002 2746
rect 17002 2694 17012 2746
rect 17036 2694 17066 2746
rect 17066 2694 17078 2746
rect 17078 2694 17092 2746
rect 17116 2694 17130 2746
rect 17130 2694 17142 2746
rect 17142 2694 17172 2746
rect 17196 2694 17206 2746
rect 17206 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 17616 2202 17672 2204
rect 17696 2202 17752 2204
rect 17776 2202 17832 2204
rect 17856 2202 17912 2204
rect 17616 2150 17662 2202
rect 17662 2150 17672 2202
rect 17696 2150 17726 2202
rect 17726 2150 17738 2202
rect 17738 2150 17752 2202
rect 17776 2150 17790 2202
rect 17790 2150 17802 2202
rect 17802 2150 17832 2202
rect 17856 2150 17866 2202
rect 17866 2150 17912 2202
rect 17616 2148 17672 2150
rect 17696 2148 17752 2150
rect 17776 2148 17832 2150
rect 17856 2148 17912 2150
rect 17866 40 17922 96
<< metal3 >>
rect 0 18458 800 18488
rect 1577 18458 1643 18461
rect 0 18456 1643 18458
rect 0 18400 1582 18456
rect 1638 18400 1643 18456
rect 0 18398 1643 18400
rect 0 18368 800 18398
rect 1577 18395 1643 18398
rect 17861 18458 17927 18461
rect 19200 18458 20000 18488
rect 17861 18456 20000 18458
rect 17861 18400 17866 18456
rect 17922 18400 20000 18456
rect 17861 18398 20000 18400
rect 17861 18395 17927 18398
rect 19200 18368 20000 18398
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 7606 17440 7922 17441
rect 7606 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7922 17440
rect 7606 17375 7922 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 17606 17440 17922 17441
rect 17606 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17922 17440
rect 17606 17375 17922 17376
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 6946 16896 7262 16897
rect 6946 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7262 16896
rect 6946 16831 7262 16832
rect 11946 16896 12262 16897
rect 11946 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12262 16896
rect 11946 16831 12262 16832
rect 16946 16896 17262 16897
rect 16946 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17262 16896
rect 16946 16831 17262 16832
rect 5349 16690 5415 16693
rect 8150 16690 8156 16692
rect 5349 16688 8156 16690
rect 5349 16632 5354 16688
rect 5410 16632 8156 16688
rect 5349 16630 8156 16632
rect 5349 16627 5415 16630
rect 8150 16628 8156 16630
rect 8220 16628 8226 16692
rect 5758 16492 5764 16556
rect 5828 16554 5834 16556
rect 13169 16554 13235 16557
rect 5828 16552 13235 16554
rect 5828 16496 13174 16552
rect 13230 16496 13235 16552
rect 5828 16494 13235 16496
rect 5828 16492 5834 16494
rect 13169 16491 13235 16494
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 7606 16352 7922 16353
rect 7606 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7922 16352
rect 7606 16287 7922 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 17606 16352 17922 16353
rect 17606 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17922 16352
rect 17606 16287 17922 16288
rect 3233 16146 3299 16149
rect 4061 16146 4127 16149
rect 12617 16146 12683 16149
rect 3233 16144 12683 16146
rect 3233 16088 3238 16144
rect 3294 16088 4066 16144
rect 4122 16088 12622 16144
rect 12678 16088 12683 16144
rect 3233 16086 12683 16088
rect 3233 16083 3299 16086
rect 4061 16083 4127 16086
rect 12617 16083 12683 16086
rect 12801 16146 12867 16149
rect 14825 16146 14891 16149
rect 12801 16144 14891 16146
rect 12801 16088 12806 16144
rect 12862 16088 14830 16144
rect 14886 16088 14891 16144
rect 12801 16086 14891 16088
rect 12801 16083 12867 16086
rect 14825 16083 14891 16086
rect 1485 16010 1551 16013
rect 7373 16010 7439 16013
rect 16389 16010 16455 16013
rect 16573 16010 16639 16013
rect 1485 16008 16639 16010
rect 1485 15952 1490 16008
rect 1546 15952 7378 16008
rect 7434 15952 16394 16008
rect 16450 15952 16578 16008
rect 16634 15952 16639 16008
rect 1485 15950 16639 15952
rect 1485 15947 1551 15950
rect 7373 15947 7439 15950
rect 16389 15947 16455 15950
rect 16573 15947 16639 15950
rect 12617 15874 12683 15877
rect 13261 15874 13327 15877
rect 12617 15872 13327 15874
rect 12617 15816 12622 15872
rect 12678 15816 13266 15872
rect 13322 15816 13327 15872
rect 12617 15814 13327 15816
rect 12617 15811 12683 15814
rect 13261 15811 13327 15814
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 16946 15808 17262 15809
rect 16946 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17262 15808
rect 16946 15743 17262 15744
rect 18229 15738 18295 15741
rect 19200 15738 20000 15768
rect 18229 15736 20000 15738
rect 18229 15680 18234 15736
rect 18290 15680 20000 15736
rect 18229 15678 20000 15680
rect 18229 15675 18295 15678
rect 19200 15648 20000 15678
rect 3969 15602 4035 15605
rect 11145 15602 11211 15605
rect 3969 15600 11211 15602
rect 3969 15544 3974 15600
rect 4030 15544 11150 15600
rect 11206 15544 11211 15600
rect 3969 15542 11211 15544
rect 3969 15539 4035 15542
rect 11145 15539 11211 15542
rect 11973 15602 12039 15605
rect 14273 15602 14339 15605
rect 11973 15600 14339 15602
rect 11973 15544 11978 15600
rect 12034 15544 14278 15600
rect 14334 15544 14339 15600
rect 11973 15542 14339 15544
rect 11973 15539 12039 15542
rect 14273 15539 14339 15542
rect 6729 15466 6795 15469
rect 14365 15466 14431 15469
rect 6729 15464 14431 15466
rect 6729 15408 6734 15464
rect 6790 15408 14370 15464
rect 14426 15408 14431 15464
rect 6729 15406 14431 15408
rect 6729 15403 6795 15406
rect 14365 15403 14431 15406
rect 5165 15330 5231 15333
rect 5390 15330 5396 15332
rect 5165 15328 5396 15330
rect 5165 15272 5170 15328
rect 5226 15272 5396 15328
rect 5165 15270 5396 15272
rect 5165 15267 5231 15270
rect 5390 15268 5396 15270
rect 5460 15268 5466 15332
rect 9121 15330 9187 15333
rect 9622 15330 9628 15332
rect 9121 15328 9628 15330
rect 9121 15272 9126 15328
rect 9182 15272 9628 15328
rect 9121 15270 9628 15272
rect 9121 15267 9187 15270
rect 9622 15268 9628 15270
rect 9692 15268 9698 15332
rect 10593 15330 10659 15333
rect 12433 15330 12499 15333
rect 13905 15332 13971 15333
rect 15009 15332 15075 15333
rect 13854 15330 13860 15332
rect 10593 15328 12499 15330
rect 10593 15272 10598 15328
rect 10654 15272 12438 15328
rect 12494 15272 12499 15328
rect 10593 15270 12499 15272
rect 13814 15270 13860 15330
rect 13924 15328 13971 15332
rect 14958 15330 14964 15332
rect 13966 15272 13971 15328
rect 10593 15267 10659 15270
rect 12433 15267 12499 15270
rect 13854 15268 13860 15270
rect 13924 15268 13971 15272
rect 14918 15270 14964 15330
rect 15028 15328 15075 15332
rect 15070 15272 15075 15328
rect 14958 15268 14964 15270
rect 15028 15268 15075 15272
rect 13905 15267 13971 15268
rect 15009 15267 15075 15268
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 17606 15264 17922 15265
rect 17606 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17922 15264
rect 17606 15199 17922 15200
rect 10777 15194 10843 15197
rect 11881 15194 11947 15197
rect 10777 15192 11947 15194
rect 10777 15136 10782 15192
rect 10838 15136 11886 15192
rect 11942 15136 11947 15192
rect 10777 15134 11947 15136
rect 10777 15131 10843 15134
rect 11881 15131 11947 15134
rect 0 15058 800 15088
rect 1577 15058 1643 15061
rect 0 15056 1643 15058
rect 0 15000 1582 15056
rect 1638 15000 1643 15056
rect 0 14998 1643 15000
rect 0 14968 800 14998
rect 1577 14995 1643 14998
rect 8661 15058 8727 15061
rect 12157 15058 12223 15061
rect 8661 15056 12223 15058
rect 8661 15000 8666 15056
rect 8722 15000 12162 15056
rect 12218 15000 12223 15056
rect 8661 14998 12223 15000
rect 8661 14995 8727 14998
rect 12157 14995 12223 14998
rect 5206 14860 5212 14924
rect 5276 14922 5282 14924
rect 16941 14922 17007 14925
rect 5276 14920 17007 14922
rect 5276 14864 16946 14920
rect 17002 14864 17007 14920
rect 5276 14862 17007 14864
rect 5276 14860 5282 14862
rect 16941 14859 17007 14862
rect 10685 14786 10751 14789
rect 11605 14786 11671 14789
rect 10685 14784 11671 14786
rect 10685 14728 10690 14784
rect 10746 14728 11610 14784
rect 11666 14728 11671 14784
rect 10685 14726 11671 14728
rect 10685 14723 10751 14726
rect 11605 14723 11671 14726
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 16946 14720 17262 14721
rect 16946 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17262 14720
rect 16946 14655 17262 14656
rect 4797 14514 4863 14517
rect 11973 14514 12039 14517
rect 4797 14512 12039 14514
rect 4797 14456 4802 14512
rect 4858 14456 11978 14512
rect 12034 14456 12039 14512
rect 4797 14454 12039 14456
rect 4797 14451 4863 14454
rect 11973 14451 12039 14454
rect 3417 14378 3483 14381
rect 11421 14378 11487 14381
rect 12893 14378 12959 14381
rect 3417 14376 11487 14378
rect 3417 14320 3422 14376
rect 3478 14320 11426 14376
rect 11482 14320 11487 14376
rect 3417 14318 11487 14320
rect 3417 14315 3483 14318
rect 11421 14315 11487 14318
rect 11608 14376 12959 14378
rect 11608 14320 12898 14376
rect 12954 14320 12959 14376
rect 11608 14318 12959 14320
rect 10317 14242 10383 14245
rect 11608 14242 11668 14318
rect 12893 14315 12959 14318
rect 10317 14240 11668 14242
rect 10317 14184 10322 14240
rect 10378 14184 11668 14240
rect 10317 14182 11668 14184
rect 10317 14179 10383 14182
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 17606 14176 17922 14177
rect 17606 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17922 14176
rect 17606 14111 17922 14112
rect 2497 13970 2563 13973
rect 6361 13970 6427 13973
rect 2497 13968 6427 13970
rect 2497 13912 2502 13968
rect 2558 13912 6366 13968
rect 6422 13912 6427 13968
rect 2497 13910 6427 13912
rect 2497 13907 2563 13910
rect 6361 13907 6427 13910
rect 4061 13836 4127 13837
rect 4061 13832 4108 13836
rect 4172 13834 4178 13836
rect 4337 13834 4403 13837
rect 8201 13834 8267 13837
rect 4061 13776 4066 13832
rect 4061 13772 4108 13776
rect 4172 13774 4218 13834
rect 4337 13832 8267 13834
rect 4337 13776 4342 13832
rect 4398 13776 8206 13832
rect 8262 13776 8267 13832
rect 4337 13774 8267 13776
rect 4172 13772 4178 13774
rect 4061 13771 4127 13772
rect 4337 13771 4403 13774
rect 8201 13771 8267 13774
rect 8886 13772 8892 13836
rect 8956 13834 8962 13836
rect 15285 13834 15351 13837
rect 8956 13832 15351 13834
rect 8956 13776 15290 13832
rect 15346 13776 15351 13832
rect 8956 13774 15351 13776
rect 8956 13772 8962 13774
rect 15285 13771 15351 13774
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 16946 13632 17262 13633
rect 16946 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17262 13632
rect 16946 13567 17262 13568
rect 5165 13426 5231 13429
rect 16757 13426 16823 13429
rect 5165 13424 16823 13426
rect 5165 13368 5170 13424
rect 5226 13368 16762 13424
rect 16818 13368 16823 13424
rect 5165 13366 16823 13368
rect 5165 13363 5231 13366
rect 16757 13363 16823 13366
rect 3182 13228 3188 13292
rect 3252 13290 3258 13292
rect 13813 13290 13879 13293
rect 3252 13288 13879 13290
rect 3252 13232 13818 13288
rect 13874 13232 13879 13288
rect 3252 13230 13879 13232
rect 3252 13228 3258 13230
rect 13813 13227 13879 13230
rect 15694 13092 15700 13156
rect 15764 13154 15770 13156
rect 16297 13154 16363 13157
rect 15764 13152 16363 13154
rect 15764 13096 16302 13152
rect 16358 13096 16363 13152
rect 15764 13094 16363 13096
rect 15764 13092 15770 13094
rect 16297 13091 16363 13094
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 17606 13088 17922 13089
rect 17606 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17922 13088
rect 17606 13023 17922 13024
rect 2129 12882 2195 12885
rect 5022 12882 5028 12884
rect 2129 12880 5028 12882
rect 2129 12824 2134 12880
rect 2190 12824 5028 12880
rect 2129 12822 5028 12824
rect 2129 12819 2195 12822
rect 5022 12820 5028 12822
rect 5092 12820 5098 12884
rect 6361 12882 6427 12885
rect 12249 12882 12315 12885
rect 6361 12880 12315 12882
rect 6361 12824 6366 12880
rect 6422 12824 12254 12880
rect 12310 12824 12315 12880
rect 6361 12822 12315 12824
rect 6361 12819 6427 12822
rect 12249 12819 12315 12822
rect 4521 12746 4587 12749
rect 12985 12746 13051 12749
rect 16849 12748 16915 12749
rect 16798 12746 16804 12748
rect 4521 12744 13051 12746
rect 4521 12688 4526 12744
rect 4582 12688 12990 12744
rect 13046 12688 13051 12744
rect 4521 12686 13051 12688
rect 16758 12686 16804 12746
rect 16868 12744 16915 12748
rect 16910 12688 16915 12744
rect 4521 12683 4587 12686
rect 12985 12683 13051 12686
rect 16798 12684 16804 12686
rect 16868 12684 16915 12688
rect 16849 12683 16915 12684
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 16946 12544 17262 12545
rect 16946 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17262 12544
rect 16946 12479 17262 12480
rect 7741 12474 7807 12477
rect 8334 12474 8340 12476
rect 7741 12472 8340 12474
rect 7741 12416 7746 12472
rect 7802 12416 8340 12472
rect 7741 12414 8340 12416
rect 7741 12411 7807 12414
rect 8334 12412 8340 12414
rect 8404 12412 8410 12476
rect 0 12338 800 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 3049 12338 3115 12341
rect 8477 12338 8543 12341
rect 3049 12336 8543 12338
rect 3049 12280 3054 12336
rect 3110 12280 8482 12336
rect 8538 12280 8543 12336
rect 3049 12278 8543 12280
rect 3049 12275 3115 12278
rect 8477 12275 8543 12278
rect 10225 12338 10291 12341
rect 14917 12338 14983 12341
rect 16757 12340 16823 12341
rect 16757 12338 16804 12340
rect 10225 12336 14983 12338
rect 10225 12280 10230 12336
rect 10286 12280 14922 12336
rect 14978 12280 14983 12336
rect 10225 12278 14983 12280
rect 16712 12336 16804 12338
rect 16712 12280 16762 12336
rect 16712 12278 16804 12280
rect 10225 12275 10291 12278
rect 14917 12275 14983 12278
rect 16757 12276 16804 12278
rect 16868 12276 16874 12340
rect 18137 12338 18203 12341
rect 19200 12338 20000 12368
rect 18137 12336 20000 12338
rect 18137 12280 18142 12336
rect 18198 12280 20000 12336
rect 18137 12278 20000 12280
rect 16757 12275 16823 12276
rect 18137 12275 18203 12278
rect 19200 12248 20000 12278
rect 2865 12202 2931 12205
rect 4153 12202 4219 12205
rect 2865 12200 4219 12202
rect 2865 12144 2870 12200
rect 2926 12144 4158 12200
rect 4214 12144 4219 12200
rect 2865 12142 4219 12144
rect 2865 12139 2931 12142
rect 4153 12139 4219 12142
rect 5349 12202 5415 12205
rect 14089 12202 14155 12205
rect 5349 12200 14155 12202
rect 5349 12144 5354 12200
rect 5410 12144 14094 12200
rect 14150 12144 14155 12200
rect 5349 12142 14155 12144
rect 5349 12139 5415 12142
rect 14089 12139 14155 12142
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 17606 12000 17922 12001
rect 17606 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17922 12000
rect 17606 11935 17922 11936
rect 7414 11930 7420 11932
rect 5950 11870 7420 11930
rect 1945 11794 2011 11797
rect 2221 11794 2287 11797
rect 5950 11794 6010 11870
rect 7414 11868 7420 11870
rect 7484 11868 7490 11932
rect 10041 11930 10107 11933
rect 11881 11930 11947 11933
rect 10041 11928 11947 11930
rect 10041 11872 10046 11928
rect 10102 11872 11886 11928
rect 11942 11872 11947 11928
rect 10041 11870 11947 11872
rect 10041 11867 10107 11870
rect 11881 11867 11947 11870
rect 1945 11792 6010 11794
rect 1945 11736 1950 11792
rect 2006 11736 2226 11792
rect 2282 11736 6010 11792
rect 1945 11734 6010 11736
rect 6085 11794 6151 11797
rect 15101 11794 15167 11797
rect 6085 11792 15167 11794
rect 6085 11736 6090 11792
rect 6146 11736 15106 11792
rect 15162 11736 15167 11792
rect 6085 11734 15167 11736
rect 1945 11731 2011 11734
rect 2221 11731 2287 11734
rect 6085 11731 6151 11734
rect 15101 11731 15167 11734
rect 6545 11658 6611 11661
rect 7649 11658 7715 11661
rect 6545 11656 7715 11658
rect 6545 11600 6550 11656
rect 6606 11600 7654 11656
rect 7710 11600 7715 11656
rect 6545 11598 7715 11600
rect 6545 11595 6611 11598
rect 7649 11595 7715 11598
rect 8109 11658 8175 11661
rect 13353 11658 13419 11661
rect 8109 11656 13419 11658
rect 8109 11600 8114 11656
rect 8170 11600 13358 11656
rect 13414 11600 13419 11656
rect 8109 11598 13419 11600
rect 8109 11595 8175 11598
rect 13353 11595 13419 11598
rect 9765 11524 9831 11525
rect 7414 11460 7420 11524
rect 7484 11522 7490 11524
rect 9765 11522 9812 11524
rect 7484 11520 9812 11522
rect 9876 11522 9882 11524
rect 10593 11522 10659 11525
rect 7484 11464 9770 11520
rect 7484 11462 9812 11464
rect 7484 11460 7490 11462
rect 9765 11460 9812 11462
rect 9876 11462 9958 11522
rect 10182 11520 10659 11522
rect 10182 11464 10598 11520
rect 10654 11464 10659 11520
rect 10182 11462 10659 11464
rect 9876 11460 9882 11462
rect 9765 11459 9831 11460
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 9673 11386 9739 11389
rect 10182 11388 10242 11462
rect 10593 11459 10659 11462
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 16946 11456 17262 11457
rect 16946 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17262 11456
rect 16946 11391 17262 11392
rect 10174 11386 10180 11388
rect 9673 11384 10180 11386
rect 9673 11328 9678 11384
rect 9734 11328 10180 11384
rect 9673 11326 10180 11328
rect 9673 11323 9739 11326
rect 10174 11324 10180 11326
rect 10244 11324 10250 11388
rect 10409 11386 10475 11389
rect 11053 11386 11119 11389
rect 10409 11384 11119 11386
rect 10409 11328 10414 11384
rect 10470 11328 11058 11384
rect 11114 11328 11119 11384
rect 10409 11326 11119 11328
rect 10409 11323 10475 11326
rect 11053 11323 11119 11326
rect 1761 11250 1827 11253
rect 11053 11250 11119 11253
rect 1761 11248 11119 11250
rect 1761 11192 1766 11248
rect 1822 11192 11058 11248
rect 11114 11192 11119 11248
rect 1761 11190 11119 11192
rect 1761 11187 1827 11190
rect 11053 11187 11119 11190
rect 12249 11250 12315 11253
rect 17125 11250 17191 11253
rect 12249 11248 17191 11250
rect 12249 11192 12254 11248
rect 12310 11192 17130 11248
rect 17186 11192 17191 11248
rect 12249 11190 17191 11192
rect 12249 11187 12315 11190
rect 17125 11187 17191 11190
rect 3877 11114 3943 11117
rect 8845 11114 8911 11117
rect 3877 11112 8911 11114
rect 3877 11056 3882 11112
rect 3938 11056 8850 11112
rect 8906 11056 8911 11112
rect 3877 11054 8911 11056
rect 3877 11051 3943 11054
rect 8845 11051 8911 11054
rect 9121 11114 9187 11117
rect 9438 11114 9444 11116
rect 9121 11112 9444 11114
rect 9121 11056 9126 11112
rect 9182 11056 9444 11112
rect 9121 11054 9444 11056
rect 9121 11051 9187 11054
rect 9438 11052 9444 11054
rect 9508 11052 9514 11116
rect 10225 11114 10291 11117
rect 10961 11114 11027 11117
rect 10225 11112 11027 11114
rect 10225 11056 10230 11112
rect 10286 11056 10966 11112
rect 11022 11056 11027 11112
rect 10225 11054 11027 11056
rect 10225 11051 10291 11054
rect 10961 11051 11027 11054
rect 5073 10978 5139 10981
rect 10225 10980 10291 10981
rect 6678 10978 6684 10980
rect 5073 10976 6684 10978
rect 5073 10920 5078 10976
rect 5134 10920 6684 10976
rect 5073 10918 6684 10920
rect 5073 10915 5139 10918
rect 6678 10916 6684 10918
rect 6748 10916 6754 10980
rect 10174 10978 10180 10980
rect 10134 10918 10180 10978
rect 10244 10976 10291 10980
rect 10286 10920 10291 10976
rect 10174 10916 10180 10918
rect 10244 10916 10291 10920
rect 10225 10915 10291 10916
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 17606 10912 17922 10913
rect 17606 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17922 10912
rect 17606 10847 17922 10848
rect 15469 10842 15535 10845
rect 15837 10842 15903 10845
rect 15469 10840 15903 10842
rect 15469 10784 15474 10840
rect 15530 10784 15842 10840
rect 15898 10784 15903 10840
rect 15469 10782 15903 10784
rect 15469 10779 15535 10782
rect 15837 10779 15903 10782
rect 4429 10706 4495 10709
rect 8477 10706 8543 10709
rect 4429 10704 8543 10706
rect 4429 10648 4434 10704
rect 4490 10648 8482 10704
rect 8538 10648 8543 10704
rect 4429 10646 8543 10648
rect 4429 10643 4495 10646
rect 8477 10643 8543 10646
rect 9622 10644 9628 10708
rect 9692 10706 9698 10708
rect 13353 10706 13419 10709
rect 9692 10704 13419 10706
rect 9692 10648 13358 10704
rect 13414 10648 13419 10704
rect 9692 10646 13419 10648
rect 9692 10644 9698 10646
rect 13353 10643 13419 10646
rect 2497 10570 2563 10573
rect 11094 10570 11100 10572
rect 2497 10568 11100 10570
rect 2497 10512 2502 10568
rect 2558 10512 11100 10568
rect 2497 10510 11100 10512
rect 2497 10507 2563 10510
rect 11094 10508 11100 10510
rect 11164 10508 11170 10572
rect 13629 10570 13695 10573
rect 13629 10568 13738 10570
rect 13629 10512 13634 10568
rect 13690 10512 13738 10568
rect 13629 10507 13738 10512
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 13678 10301 13738 10507
rect 16946 10368 17262 10369
rect 16946 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17262 10368
rect 16946 10303 17262 10304
rect 2497 10298 2563 10301
rect 5257 10298 5323 10301
rect 2497 10296 5323 10298
rect 2497 10240 2502 10296
rect 2558 10240 5262 10296
rect 5318 10240 5323 10296
rect 2497 10238 5323 10240
rect 2497 10235 2563 10238
rect 5257 10235 5323 10238
rect 13629 10296 13738 10301
rect 13629 10240 13634 10296
rect 13690 10240 13738 10296
rect 13629 10238 13738 10240
rect 13629 10235 13695 10238
rect 11237 10162 11303 10165
rect 12525 10162 12591 10165
rect 11237 10160 12591 10162
rect 11237 10104 11242 10160
rect 11298 10104 12530 10160
rect 12586 10104 12591 10160
rect 11237 10102 12591 10104
rect 11237 10099 11303 10102
rect 12525 10099 12591 10102
rect 3049 10026 3115 10029
rect 8569 10026 8635 10029
rect 3049 10024 8635 10026
rect 3049 9968 3054 10024
rect 3110 9968 8574 10024
rect 8630 9968 8635 10024
rect 3049 9966 8635 9968
rect 3049 9963 3115 9966
rect 8569 9963 8635 9966
rect 8293 9892 8359 9893
rect 8293 9890 8340 9892
rect 8248 9888 8340 9890
rect 8248 9832 8298 9888
rect 8248 9830 8340 9832
rect 8293 9828 8340 9830
rect 8404 9828 8410 9892
rect 8293 9827 8359 9828
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 17606 9824 17922 9825
rect 17606 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17922 9824
rect 17606 9759 17922 9760
rect 7189 9754 7255 9757
rect 7414 9754 7420 9756
rect 7189 9752 7420 9754
rect 7189 9696 7194 9752
rect 7250 9696 7420 9752
rect 7189 9694 7420 9696
rect 7189 9691 7255 9694
rect 7414 9692 7420 9694
rect 7484 9692 7490 9756
rect 8661 9754 8727 9757
rect 8112 9752 8727 9754
rect 8112 9696 8666 9752
rect 8722 9696 8727 9752
rect 8112 9694 8727 9696
rect 8112 9652 8172 9694
rect 8661 9691 8727 9694
rect 15142 9692 15148 9756
rect 15212 9754 15218 9756
rect 15377 9754 15443 9757
rect 15212 9752 15443 9754
rect 15212 9696 15382 9752
rect 15438 9696 15443 9752
rect 15212 9694 15443 9696
rect 15212 9692 15218 9694
rect 15377 9691 15443 9694
rect 7974 9621 8172 9652
rect 5022 9556 5028 9620
rect 5092 9618 5098 9620
rect 5165 9618 5231 9621
rect 5092 9616 5231 9618
rect 5092 9560 5170 9616
rect 5226 9560 5231 9616
rect 5092 9558 5231 9560
rect 5092 9556 5098 9558
rect 5165 9555 5231 9558
rect 7925 9616 8172 9621
rect 17401 9618 17467 9621
rect 7925 9560 7930 9616
rect 7986 9592 8172 9616
rect 8250 9616 17467 9618
rect 7986 9560 8034 9592
rect 7925 9558 8034 9560
rect 8250 9560 17406 9616
rect 17462 9560 17467 9616
rect 8250 9558 17467 9560
rect 7925 9555 7991 9558
rect 6085 9482 6151 9485
rect 6913 9482 6979 9485
rect 6085 9480 6979 9482
rect 6085 9424 6090 9480
rect 6146 9424 6918 9480
rect 6974 9424 6979 9480
rect 6085 9422 6979 9424
rect 6085 9419 6151 9422
rect 6913 9419 6979 9422
rect 7465 9346 7531 9349
rect 8250 9346 8310 9558
rect 17401 9555 17467 9558
rect 18137 9618 18203 9621
rect 19200 9618 20000 9648
rect 18137 9616 20000 9618
rect 18137 9560 18142 9616
rect 18198 9560 20000 9616
rect 18137 9558 20000 9560
rect 18137 9555 18203 9558
rect 19200 9528 20000 9558
rect 10501 9482 10567 9485
rect 12433 9482 12499 9485
rect 10501 9480 12499 9482
rect 10501 9424 10506 9480
rect 10562 9424 12438 9480
rect 12494 9424 12499 9480
rect 10501 9422 12499 9424
rect 10501 9419 10567 9422
rect 12433 9419 12499 9422
rect 7465 9344 8310 9346
rect 7465 9288 7470 9344
rect 7526 9288 8310 9344
rect 7465 9286 8310 9288
rect 7465 9283 7531 9286
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 16946 9280 17262 9281
rect 16946 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17262 9280
rect 16946 9215 17262 9216
rect 7465 9212 7531 9213
rect 7414 9148 7420 9212
rect 7484 9210 7531 9212
rect 7484 9208 7576 9210
rect 7526 9152 7576 9208
rect 7484 9150 7576 9152
rect 7484 9148 7531 9150
rect 7465 9147 7531 9148
rect 5533 9074 5599 9077
rect 13854 9074 13860 9076
rect 5533 9072 13860 9074
rect 5533 9016 5538 9072
rect 5594 9016 13860 9072
rect 5533 9014 13860 9016
rect 5533 9011 5599 9014
rect 13854 9012 13860 9014
rect 13924 9012 13930 9076
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 17606 8736 17922 8737
rect 17606 8672 17612 8736
rect 17676 8672 17692 8736
rect 17756 8672 17772 8736
rect 17836 8672 17852 8736
rect 17916 8672 17922 8736
rect 17606 8671 17922 8672
rect 8201 8668 8267 8669
rect 8150 8604 8156 8668
rect 8220 8666 8267 8668
rect 8220 8664 8312 8666
rect 8262 8608 8312 8664
rect 8220 8606 8312 8608
rect 8220 8604 8267 8606
rect 8201 8603 8267 8604
rect 5717 8530 5783 8533
rect 9397 8530 9463 8533
rect 5717 8528 9463 8530
rect 5717 8472 5722 8528
rect 5778 8472 9402 8528
rect 9458 8472 9463 8528
rect 5717 8470 9463 8472
rect 5717 8467 5783 8470
rect 9397 8467 9463 8470
rect 13445 8530 13511 8533
rect 13813 8530 13879 8533
rect 13445 8528 13879 8530
rect 13445 8472 13450 8528
rect 13506 8472 13818 8528
rect 13874 8472 13879 8528
rect 13445 8470 13879 8472
rect 13445 8467 13511 8470
rect 13813 8467 13879 8470
rect 9806 8332 9812 8396
rect 9876 8394 9882 8396
rect 9876 8334 13554 8394
rect 9876 8332 9882 8334
rect 13494 8261 13554 8334
rect 13494 8256 13603 8261
rect 13494 8200 13542 8256
rect 13598 8200 13603 8256
rect 13494 8198 13603 8200
rect 13537 8195 13603 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 16946 8192 17262 8193
rect 16946 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17262 8192
rect 16946 8127 17262 8128
rect 9857 8122 9923 8125
rect 8158 8120 9923 8122
rect 8158 8064 9862 8120
rect 9918 8064 9923 8120
rect 8158 8062 9923 8064
rect 3693 7986 3759 7989
rect 8158 7986 8218 8062
rect 9857 8059 9923 8062
rect 3693 7984 8218 7986
rect 3693 7928 3698 7984
rect 3754 7928 8218 7984
rect 3693 7926 8218 7928
rect 8385 7986 8451 7989
rect 15142 7986 15148 7988
rect 8385 7984 15148 7986
rect 8385 7928 8390 7984
rect 8446 7928 15148 7984
rect 8385 7926 15148 7928
rect 3693 7923 3759 7926
rect 8385 7923 8451 7926
rect 15142 7924 15148 7926
rect 15212 7924 15218 7988
rect 6494 7788 6500 7852
rect 6564 7850 6570 7852
rect 7097 7850 7163 7853
rect 6564 7848 7163 7850
rect 6564 7792 7102 7848
rect 7158 7792 7163 7848
rect 6564 7790 7163 7792
rect 6564 7788 6570 7790
rect 7097 7787 7163 7790
rect 7281 7850 7347 7853
rect 18321 7850 18387 7853
rect 7281 7848 18387 7850
rect 7281 7792 7286 7848
rect 7342 7792 18326 7848
rect 18382 7792 18387 7848
rect 7281 7790 18387 7792
rect 7281 7787 7347 7790
rect 18321 7787 18387 7790
rect 5993 7714 6059 7717
rect 6545 7714 6611 7717
rect 6729 7714 6795 7717
rect 5993 7712 6795 7714
rect 5993 7656 5998 7712
rect 6054 7656 6550 7712
rect 6606 7656 6734 7712
rect 6790 7656 6795 7712
rect 5993 7654 6795 7656
rect 5993 7651 6059 7654
rect 6545 7651 6611 7654
rect 6729 7651 6795 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 17606 7648 17922 7649
rect 17606 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17922 7648
rect 17606 7583 17922 7584
rect 6269 7578 6335 7581
rect 6913 7578 6979 7581
rect 6269 7576 6979 7578
rect 6269 7520 6274 7576
rect 6330 7520 6918 7576
rect 6974 7520 6979 7576
rect 6269 7518 6979 7520
rect 6269 7515 6335 7518
rect 6913 7515 6979 7518
rect 4102 7380 4108 7444
rect 4172 7442 4178 7444
rect 16389 7442 16455 7445
rect 4172 7440 16455 7442
rect 4172 7384 16394 7440
rect 16450 7384 16455 7440
rect 4172 7382 16455 7384
rect 4172 7380 4178 7382
rect 16389 7379 16455 7382
rect 3693 7306 3759 7309
rect 8201 7306 8267 7309
rect 3693 7304 8267 7306
rect 3693 7248 3698 7304
rect 3754 7248 8206 7304
rect 8262 7248 8267 7304
rect 3693 7246 8267 7248
rect 3693 7243 3759 7246
rect 8201 7243 8267 7246
rect 5717 7170 5783 7173
rect 6729 7172 6795 7173
rect 6494 7170 6500 7172
rect 5717 7168 6500 7170
rect 5717 7112 5722 7168
rect 5778 7112 6500 7168
rect 5717 7110 6500 7112
rect 5717 7107 5783 7110
rect 6494 7108 6500 7110
rect 6564 7108 6570 7172
rect 6678 7108 6684 7172
rect 6748 7170 6795 7172
rect 6748 7168 6840 7170
rect 6790 7112 6840 7168
rect 6748 7110 6840 7112
rect 6748 7108 6795 7110
rect 6729 7107 6795 7108
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 16946 7104 17262 7105
rect 16946 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17262 7104
rect 16946 7039 17262 7040
rect 5390 6972 5396 7036
rect 5460 7034 5466 7036
rect 6545 7034 6611 7037
rect 5460 7032 6611 7034
rect 5460 6976 6550 7032
rect 6606 6976 6611 7032
rect 5460 6974 6611 6976
rect 5460 6972 5466 6974
rect 6545 6971 6611 6974
rect 3785 6898 3851 6901
rect 5717 6900 5783 6901
rect 3785 6896 5642 6898
rect 3785 6840 3790 6896
rect 3846 6840 5642 6896
rect 3785 6838 5642 6840
rect 3785 6835 3851 6838
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 0 6218 800 6248
rect 933 6218 999 6221
rect 0 6216 999 6218
rect 0 6160 938 6216
rect 994 6160 999 6216
rect 0 6158 999 6160
rect 0 6128 800 6158
rect 933 6155 999 6158
rect 1945 6218 2011 6221
rect 5582 6218 5642 6838
rect 5717 6896 5764 6900
rect 5828 6898 5834 6900
rect 6729 6898 6795 6901
rect 14641 6898 14707 6901
rect 5717 6840 5722 6896
rect 5717 6836 5764 6840
rect 5828 6838 5874 6898
rect 6729 6896 14707 6898
rect 6729 6840 6734 6896
rect 6790 6840 14646 6896
rect 14702 6840 14707 6896
rect 6729 6838 14707 6840
rect 5828 6836 5834 6838
rect 5717 6835 5783 6836
rect 6729 6835 6795 6838
rect 11654 6765 11714 6838
rect 14641 6835 14707 6838
rect 5809 6762 5875 6765
rect 11053 6762 11119 6765
rect 5809 6760 11119 6762
rect 5809 6704 5814 6760
rect 5870 6704 11058 6760
rect 11114 6704 11119 6760
rect 5809 6702 11119 6704
rect 11654 6760 11763 6765
rect 15377 6762 15443 6765
rect 11654 6704 11702 6760
rect 11758 6704 11763 6760
rect 11654 6702 11763 6704
rect 5809 6699 5875 6702
rect 11053 6699 11119 6702
rect 11697 6699 11763 6702
rect 12390 6760 15443 6762
rect 12390 6704 15382 6760
rect 15438 6704 15443 6760
rect 12390 6702 15443 6704
rect 8753 6626 8819 6629
rect 12390 6626 12450 6702
rect 15377 6699 15443 6702
rect 8753 6624 12450 6626
rect 8753 6568 8758 6624
rect 8814 6568 12450 6624
rect 8753 6566 12450 6568
rect 8753 6563 8819 6566
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 17606 6560 17922 6561
rect 17606 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17922 6560
rect 17606 6495 17922 6496
rect 11421 6490 11487 6493
rect 11605 6490 11671 6493
rect 11421 6488 11671 6490
rect 11421 6432 11426 6488
rect 11482 6432 11610 6488
rect 11666 6432 11671 6488
rect 11421 6430 11671 6432
rect 11421 6427 11487 6430
rect 11605 6427 11671 6430
rect 6637 6354 6703 6357
rect 17953 6354 18019 6357
rect 6637 6352 18019 6354
rect 6637 6296 6642 6352
rect 6698 6296 17958 6352
rect 18014 6296 18019 6352
rect 6637 6294 18019 6296
rect 6637 6291 6703 6294
rect 17953 6291 18019 6294
rect 8293 6218 8359 6221
rect 13813 6218 13879 6221
rect 1945 6216 2514 6218
rect 1945 6160 1950 6216
rect 2006 6160 2514 6216
rect 1945 6158 2514 6160
rect 5582 6158 8218 6218
rect 1945 6155 2011 6158
rect 2454 6082 2514 6158
rect 5625 6082 5691 6085
rect 6637 6082 6703 6085
rect 2454 6080 6703 6082
rect 2454 6024 5630 6080
rect 5686 6024 6642 6080
rect 6698 6024 6703 6080
rect 2454 6022 6703 6024
rect 8158 6082 8218 6158
rect 8293 6216 13879 6218
rect 8293 6160 8298 6216
rect 8354 6160 13818 6216
rect 13874 6160 13879 6216
rect 8293 6158 13879 6160
rect 8293 6155 8359 6158
rect 13813 6155 13879 6158
rect 18413 6218 18479 6221
rect 19200 6218 20000 6248
rect 18413 6216 20000 6218
rect 18413 6160 18418 6216
rect 18474 6160 20000 6216
rect 18413 6158 20000 6160
rect 18413 6155 18479 6158
rect 19200 6128 20000 6158
rect 8753 6082 8819 6085
rect 8158 6080 8819 6082
rect 8158 6024 8758 6080
rect 8814 6024 8819 6080
rect 8158 6022 8819 6024
rect 5625 6019 5691 6022
rect 6637 6019 6703 6022
rect 8753 6019 8819 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 16946 6016 17262 6017
rect 16946 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17262 6016
rect 16946 5951 17262 5952
rect 7833 5946 7899 5949
rect 8661 5946 8727 5949
rect 7833 5944 8727 5946
rect 7833 5888 7838 5944
rect 7894 5888 8666 5944
rect 8722 5888 8727 5944
rect 7833 5886 8727 5888
rect 7833 5883 7899 5886
rect 8661 5883 8727 5886
rect 6821 5810 6887 5813
rect 8886 5810 8892 5812
rect 6821 5808 8892 5810
rect 6821 5752 6826 5808
rect 6882 5752 8892 5808
rect 6821 5750 8892 5752
rect 6821 5747 6887 5750
rect 8886 5748 8892 5750
rect 8956 5748 8962 5812
rect 1577 5674 1643 5677
rect 14958 5674 14964 5676
rect 1577 5672 14964 5674
rect 1577 5616 1582 5672
rect 1638 5616 14964 5672
rect 1577 5614 14964 5616
rect 1577 5611 1643 5614
rect 14958 5612 14964 5614
rect 15028 5612 15034 5676
rect 3049 5538 3115 5541
rect 3182 5538 3188 5540
rect 3049 5536 3188 5538
rect 3049 5480 3054 5536
rect 3110 5480 3188 5536
rect 3049 5478 3188 5480
rect 3049 5475 3115 5478
rect 3182 5476 3188 5478
rect 3252 5476 3258 5540
rect 3601 5538 3667 5541
rect 4245 5538 4311 5541
rect 3601 5536 4311 5538
rect 3601 5480 3606 5536
rect 3662 5480 4250 5536
rect 4306 5480 4311 5536
rect 3601 5478 4311 5480
rect 3601 5475 3667 5478
rect 4245 5475 4311 5478
rect 6085 5538 6151 5541
rect 6678 5538 6684 5540
rect 6085 5536 6684 5538
rect 6085 5480 6090 5536
rect 6146 5480 6684 5536
rect 6085 5478 6684 5480
rect 6085 5475 6151 5478
rect 6678 5476 6684 5478
rect 6748 5476 6754 5540
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 17606 5472 17922 5473
rect 17606 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17922 5472
rect 17606 5407 17922 5408
rect 2405 5266 2471 5269
rect 7649 5266 7715 5269
rect 16757 5266 16823 5269
rect 2405 5264 7482 5266
rect 2405 5208 2410 5264
rect 2466 5208 7482 5264
rect 2405 5206 7482 5208
rect 2405 5203 2471 5206
rect 2037 5130 2103 5133
rect 4981 5130 5047 5133
rect 2037 5128 5047 5130
rect 2037 5072 2042 5128
rect 2098 5072 4986 5128
rect 5042 5072 5047 5128
rect 2037 5070 5047 5072
rect 7422 5130 7482 5206
rect 7649 5264 16823 5266
rect 7649 5208 7654 5264
rect 7710 5208 16762 5264
rect 16818 5208 16823 5264
rect 7649 5206 16823 5208
rect 7649 5203 7715 5206
rect 16757 5203 16823 5206
rect 9397 5130 9463 5133
rect 7422 5128 9463 5130
rect 7422 5072 9402 5128
rect 9458 5072 9463 5128
rect 7422 5070 9463 5072
rect 2037 5067 2103 5070
rect 4981 5067 5047 5070
rect 9397 5067 9463 5070
rect 10869 5130 10935 5133
rect 13721 5130 13787 5133
rect 10869 5128 13787 5130
rect 10869 5072 10874 5128
rect 10930 5072 13726 5128
rect 13782 5072 13787 5128
rect 10869 5070 13787 5072
rect 10869 5067 10935 5070
rect 13721 5067 13787 5070
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 16946 4928 17262 4929
rect 16946 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17262 4928
rect 16946 4863 17262 4864
rect 5257 4860 5323 4861
rect 5206 4796 5212 4860
rect 5276 4858 5323 4860
rect 7649 4858 7715 4861
rect 11421 4858 11487 4861
rect 5276 4856 5368 4858
rect 5318 4800 5368 4856
rect 5276 4798 5368 4800
rect 7649 4856 11487 4858
rect 7649 4800 7654 4856
rect 7710 4800 11426 4856
rect 11482 4800 11487 4856
rect 7649 4798 11487 4800
rect 5276 4796 5323 4798
rect 5257 4795 5323 4796
rect 7649 4795 7715 4798
rect 11421 4795 11487 4798
rect 4245 4722 4311 4725
rect 8201 4722 8267 4725
rect 4245 4720 8267 4722
rect 4245 4664 4250 4720
rect 4306 4664 8206 4720
rect 8262 4664 8267 4720
rect 4245 4662 8267 4664
rect 4245 4659 4311 4662
rect 8201 4659 8267 4662
rect 9673 4722 9739 4725
rect 11881 4722 11947 4725
rect 9673 4720 11947 4722
rect 9673 4664 9678 4720
rect 9734 4664 11886 4720
rect 11942 4664 11947 4720
rect 9673 4662 11947 4664
rect 9673 4659 9739 4662
rect 11881 4659 11947 4662
rect 6085 4586 6151 4589
rect 9949 4586 10015 4589
rect 10133 4586 10199 4589
rect 6085 4584 10199 4586
rect 6085 4528 6090 4584
rect 6146 4528 9954 4584
rect 10010 4528 10138 4584
rect 10194 4528 10199 4584
rect 6085 4526 10199 4528
rect 6085 4523 6151 4526
rect 9949 4523 10015 4526
rect 10133 4523 10199 4526
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 17606 4384 17922 4385
rect 17606 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17922 4384
rect 17606 4319 17922 4320
rect 2129 4178 2195 4181
rect 9305 4178 9371 4181
rect 2129 4176 9371 4178
rect 2129 4120 2134 4176
rect 2190 4120 9310 4176
rect 9366 4120 9371 4176
rect 2129 4118 9371 4120
rect 2129 4115 2195 4118
rect 9305 4115 9371 4118
rect 4337 4042 4403 4045
rect 10777 4042 10843 4045
rect 17493 4042 17559 4045
rect 4337 4040 10610 4042
rect 4337 3984 4342 4040
rect 4398 3984 10610 4040
rect 4337 3982 10610 3984
rect 4337 3979 4403 3982
rect 10550 3906 10610 3982
rect 10777 4040 17559 4042
rect 10777 3984 10782 4040
rect 10838 3984 17498 4040
rect 17554 3984 17559 4040
rect 10777 3982 17559 3984
rect 10777 3979 10843 3982
rect 17493 3979 17559 3982
rect 11789 3906 11855 3909
rect 10550 3904 11855 3906
rect 10550 3848 11794 3904
rect 11850 3848 11855 3904
rect 10550 3846 11855 3848
rect 11789 3843 11855 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 16946 3840 17262 3841
rect 16946 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17262 3840
rect 16946 3775 17262 3776
rect 11145 3772 11211 3773
rect 11094 3770 11100 3772
rect 11054 3710 11100 3770
rect 11164 3768 11211 3772
rect 11206 3712 11211 3768
rect 11094 3708 11100 3710
rect 11164 3708 11211 3712
rect 11145 3707 11211 3708
rect 9581 3634 9647 3637
rect 9581 3632 12082 3634
rect 9581 3576 9586 3632
rect 9642 3576 12082 3632
rect 9581 3574 12082 3576
rect 9581 3571 9647 3574
rect 1393 3498 1459 3501
rect 11881 3498 11947 3501
rect 1393 3496 11947 3498
rect 1393 3440 1398 3496
rect 1454 3440 11886 3496
rect 11942 3440 11947 3496
rect 1393 3438 11947 3440
rect 12022 3498 12082 3574
rect 15745 3498 15811 3501
rect 12022 3496 15811 3498
rect 12022 3440 15750 3496
rect 15806 3440 15811 3496
rect 12022 3438 15811 3440
rect 1393 3435 1459 3438
rect 11881 3435 11947 3438
rect 15745 3435 15811 3438
rect 18137 3498 18203 3501
rect 19200 3498 20000 3528
rect 18137 3496 20000 3498
rect 18137 3440 18142 3496
rect 18198 3440 20000 3496
rect 18137 3438 20000 3440
rect 18137 3435 18203 3438
rect 19200 3408 20000 3438
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 17606 3296 17922 3297
rect 17606 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17922 3296
rect 17606 3231 17922 3232
rect 12157 3226 12223 3229
rect 8158 3224 12223 3226
rect 8158 3168 12162 3224
rect 12218 3168 12223 3224
rect 8158 3166 12223 3168
rect 4337 3090 4403 3093
rect 5165 3090 5231 3093
rect 8158 3090 8218 3166
rect 12157 3163 12223 3166
rect 12341 3226 12407 3229
rect 12341 3224 12450 3226
rect 12341 3168 12346 3224
rect 12402 3168 12450 3224
rect 12341 3163 12450 3168
rect 4337 3088 8218 3090
rect 4337 3032 4342 3088
rect 4398 3032 5170 3088
rect 5226 3032 8218 3088
rect 4337 3030 8218 3032
rect 4337 3027 4403 3030
rect 5165 3027 5231 3030
rect 9438 3028 9444 3092
rect 9508 3090 9514 3092
rect 12065 3090 12131 3093
rect 9508 3088 12131 3090
rect 9508 3032 12070 3088
rect 12126 3032 12131 3088
rect 9508 3030 12131 3032
rect 12390 3090 12450 3163
rect 12525 3090 12591 3093
rect 12390 3088 12591 3090
rect 12390 3032 12530 3088
rect 12586 3032 12591 3088
rect 12390 3030 12591 3032
rect 9508 3028 9514 3030
rect 12065 3027 12131 3030
rect 12525 3027 12591 3030
rect 6545 2954 6611 2957
rect 8293 2954 8359 2957
rect 11789 2954 11855 2957
rect 6545 2952 11855 2954
rect 6545 2896 6550 2952
rect 6606 2896 8298 2952
rect 8354 2896 11794 2952
rect 11850 2896 11855 2952
rect 6545 2894 11855 2896
rect 6545 2891 6611 2894
rect 8293 2891 8359 2894
rect 11789 2891 11855 2894
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 16946 2752 17262 2753
rect 16946 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17262 2752
rect 16946 2687 17262 2688
rect 9121 2546 9187 2549
rect 15694 2546 15700 2548
rect 9121 2544 15700 2546
rect 9121 2488 9126 2544
rect 9182 2488 15700 2544
rect 9121 2486 15700 2488
rect 9121 2483 9187 2486
rect 15694 2484 15700 2486
rect 15764 2484 15770 2548
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 17606 2208 17922 2209
rect 17606 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17922 2208
rect 17606 2143 17922 2144
rect 17861 98 17927 101
rect 19200 98 20000 128
rect 17861 96 20000 98
rect 17861 40 17866 96
rect 17922 40 20000 96
rect 17861 38 20000 40
rect 17861 35 17927 38
rect 19200 8 20000 38
<< via3 >>
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 7612 17436 7676 17440
rect 7612 17380 7616 17436
rect 7616 17380 7672 17436
rect 7672 17380 7676 17436
rect 7612 17376 7676 17380
rect 7692 17436 7756 17440
rect 7692 17380 7696 17436
rect 7696 17380 7752 17436
rect 7752 17380 7756 17436
rect 7692 17376 7756 17380
rect 7772 17436 7836 17440
rect 7772 17380 7776 17436
rect 7776 17380 7832 17436
rect 7832 17380 7836 17436
rect 7772 17376 7836 17380
rect 7852 17436 7916 17440
rect 7852 17380 7856 17436
rect 7856 17380 7912 17436
rect 7912 17380 7916 17436
rect 7852 17376 7916 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 17612 17436 17676 17440
rect 17612 17380 17616 17436
rect 17616 17380 17672 17436
rect 17672 17380 17676 17436
rect 17612 17376 17676 17380
rect 17692 17436 17756 17440
rect 17692 17380 17696 17436
rect 17696 17380 17752 17436
rect 17752 17380 17756 17436
rect 17692 17376 17756 17380
rect 17772 17436 17836 17440
rect 17772 17380 17776 17436
rect 17776 17380 17832 17436
rect 17832 17380 17836 17436
rect 17772 17376 17836 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 6952 16892 7016 16896
rect 6952 16836 6956 16892
rect 6956 16836 7012 16892
rect 7012 16836 7016 16892
rect 6952 16832 7016 16836
rect 7032 16892 7096 16896
rect 7032 16836 7036 16892
rect 7036 16836 7092 16892
rect 7092 16836 7096 16892
rect 7032 16832 7096 16836
rect 7112 16892 7176 16896
rect 7112 16836 7116 16892
rect 7116 16836 7172 16892
rect 7172 16836 7176 16892
rect 7112 16832 7176 16836
rect 7192 16892 7256 16896
rect 7192 16836 7196 16892
rect 7196 16836 7252 16892
rect 7252 16836 7256 16892
rect 7192 16832 7256 16836
rect 11952 16892 12016 16896
rect 11952 16836 11956 16892
rect 11956 16836 12012 16892
rect 12012 16836 12016 16892
rect 11952 16832 12016 16836
rect 12032 16892 12096 16896
rect 12032 16836 12036 16892
rect 12036 16836 12092 16892
rect 12092 16836 12096 16892
rect 12032 16832 12096 16836
rect 12112 16892 12176 16896
rect 12112 16836 12116 16892
rect 12116 16836 12172 16892
rect 12172 16836 12176 16892
rect 12112 16832 12176 16836
rect 12192 16892 12256 16896
rect 12192 16836 12196 16892
rect 12196 16836 12252 16892
rect 12252 16836 12256 16892
rect 12192 16832 12256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 8156 16628 8220 16692
rect 5764 16492 5828 16556
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 7612 16348 7676 16352
rect 7612 16292 7616 16348
rect 7616 16292 7672 16348
rect 7672 16292 7676 16348
rect 7612 16288 7676 16292
rect 7692 16348 7756 16352
rect 7692 16292 7696 16348
rect 7696 16292 7752 16348
rect 7752 16292 7756 16348
rect 7692 16288 7756 16292
rect 7772 16348 7836 16352
rect 7772 16292 7776 16348
rect 7776 16292 7832 16348
rect 7832 16292 7836 16348
rect 7772 16288 7836 16292
rect 7852 16348 7916 16352
rect 7852 16292 7856 16348
rect 7856 16292 7912 16348
rect 7912 16292 7916 16348
rect 7852 16288 7916 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 17612 16348 17676 16352
rect 17612 16292 17616 16348
rect 17616 16292 17672 16348
rect 17672 16292 17676 16348
rect 17612 16288 17676 16292
rect 17692 16348 17756 16352
rect 17692 16292 17696 16348
rect 17696 16292 17752 16348
rect 17752 16292 17756 16348
rect 17692 16288 17756 16292
rect 17772 16348 17836 16352
rect 17772 16292 17776 16348
rect 17776 16292 17832 16348
rect 17832 16292 17836 16348
rect 17772 16288 17836 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 5396 15268 5460 15332
rect 9628 15268 9692 15332
rect 13860 15328 13924 15332
rect 13860 15272 13910 15328
rect 13910 15272 13924 15328
rect 13860 15268 13924 15272
rect 14964 15328 15028 15332
rect 14964 15272 15014 15328
rect 15014 15272 15028 15328
rect 14964 15268 15028 15272
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 17612 15260 17676 15264
rect 17612 15204 17616 15260
rect 17616 15204 17672 15260
rect 17672 15204 17676 15260
rect 17612 15200 17676 15204
rect 17692 15260 17756 15264
rect 17692 15204 17696 15260
rect 17696 15204 17752 15260
rect 17752 15204 17756 15260
rect 17692 15200 17756 15204
rect 17772 15260 17836 15264
rect 17772 15204 17776 15260
rect 17776 15204 17832 15260
rect 17832 15204 17836 15260
rect 17772 15200 17836 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 5212 14860 5276 14924
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 17612 14172 17676 14176
rect 17612 14116 17616 14172
rect 17616 14116 17672 14172
rect 17672 14116 17676 14172
rect 17612 14112 17676 14116
rect 17692 14172 17756 14176
rect 17692 14116 17696 14172
rect 17696 14116 17752 14172
rect 17752 14116 17756 14172
rect 17692 14112 17756 14116
rect 17772 14172 17836 14176
rect 17772 14116 17776 14172
rect 17776 14116 17832 14172
rect 17832 14116 17836 14172
rect 17772 14112 17836 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 4108 13832 4172 13836
rect 4108 13776 4122 13832
rect 4122 13776 4172 13832
rect 4108 13772 4172 13776
rect 8892 13772 8956 13836
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 3188 13228 3252 13292
rect 15700 13092 15764 13156
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 17612 13084 17676 13088
rect 17612 13028 17616 13084
rect 17616 13028 17672 13084
rect 17672 13028 17676 13084
rect 17612 13024 17676 13028
rect 17692 13084 17756 13088
rect 17692 13028 17696 13084
rect 17696 13028 17752 13084
rect 17752 13028 17756 13084
rect 17692 13024 17756 13028
rect 17772 13084 17836 13088
rect 17772 13028 17776 13084
rect 17776 13028 17832 13084
rect 17832 13028 17836 13084
rect 17772 13024 17836 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 5028 12820 5092 12884
rect 16804 12744 16868 12748
rect 16804 12688 16854 12744
rect 16854 12688 16868 12744
rect 16804 12684 16868 12688
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 8340 12412 8404 12476
rect 16804 12336 16868 12340
rect 16804 12280 16818 12336
rect 16818 12280 16868 12336
rect 16804 12276 16868 12280
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 17612 11996 17676 12000
rect 17612 11940 17616 11996
rect 17616 11940 17672 11996
rect 17672 11940 17676 11996
rect 17612 11936 17676 11940
rect 17692 11996 17756 12000
rect 17692 11940 17696 11996
rect 17696 11940 17752 11996
rect 17752 11940 17756 11996
rect 17692 11936 17756 11940
rect 17772 11996 17836 12000
rect 17772 11940 17776 11996
rect 17776 11940 17832 11996
rect 17832 11940 17836 11996
rect 17772 11936 17836 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 7420 11868 7484 11932
rect 7420 11460 7484 11524
rect 9812 11520 9876 11524
rect 9812 11464 9826 11520
rect 9826 11464 9876 11520
rect 9812 11460 9876 11464
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 10180 11324 10244 11388
rect 9444 11052 9508 11116
rect 6684 10916 6748 10980
rect 10180 10976 10244 10980
rect 10180 10920 10230 10976
rect 10230 10920 10244 10976
rect 10180 10916 10244 10920
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 17612 10908 17676 10912
rect 17612 10852 17616 10908
rect 17616 10852 17672 10908
rect 17672 10852 17676 10908
rect 17612 10848 17676 10852
rect 17692 10908 17756 10912
rect 17692 10852 17696 10908
rect 17696 10852 17752 10908
rect 17752 10852 17756 10908
rect 17692 10848 17756 10852
rect 17772 10908 17836 10912
rect 17772 10852 17776 10908
rect 17776 10852 17832 10908
rect 17832 10852 17836 10908
rect 17772 10848 17836 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 9628 10644 9692 10708
rect 11100 10508 11164 10572
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 8340 9888 8404 9892
rect 8340 9832 8354 9888
rect 8354 9832 8404 9888
rect 8340 9828 8404 9832
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 17612 9820 17676 9824
rect 17612 9764 17616 9820
rect 17616 9764 17672 9820
rect 17672 9764 17676 9820
rect 17612 9760 17676 9764
rect 17692 9820 17756 9824
rect 17692 9764 17696 9820
rect 17696 9764 17752 9820
rect 17752 9764 17756 9820
rect 17692 9760 17756 9764
rect 17772 9820 17836 9824
rect 17772 9764 17776 9820
rect 17776 9764 17832 9820
rect 17832 9764 17836 9820
rect 17772 9760 17836 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 7420 9692 7484 9756
rect 15148 9692 15212 9756
rect 5028 9556 5092 9620
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 7420 9208 7484 9212
rect 7420 9152 7470 9208
rect 7470 9152 7484 9208
rect 7420 9148 7484 9152
rect 13860 9012 13924 9076
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 17612 8732 17676 8736
rect 17612 8676 17616 8732
rect 17616 8676 17672 8732
rect 17672 8676 17676 8732
rect 17612 8672 17676 8676
rect 17692 8732 17756 8736
rect 17692 8676 17696 8732
rect 17696 8676 17752 8732
rect 17752 8676 17756 8732
rect 17692 8672 17756 8676
rect 17772 8732 17836 8736
rect 17772 8676 17776 8732
rect 17776 8676 17832 8732
rect 17832 8676 17836 8732
rect 17772 8672 17836 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 8156 8664 8220 8668
rect 8156 8608 8206 8664
rect 8206 8608 8220 8664
rect 8156 8604 8220 8608
rect 9812 8332 9876 8396
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 15148 7924 15212 7988
rect 6500 7788 6564 7852
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 17612 7644 17676 7648
rect 17612 7588 17616 7644
rect 17616 7588 17672 7644
rect 17672 7588 17676 7644
rect 17612 7584 17676 7588
rect 17692 7644 17756 7648
rect 17692 7588 17696 7644
rect 17696 7588 17752 7644
rect 17752 7588 17756 7644
rect 17692 7584 17756 7588
rect 17772 7644 17836 7648
rect 17772 7588 17776 7644
rect 17776 7588 17832 7644
rect 17832 7588 17836 7644
rect 17772 7584 17836 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 4108 7380 4172 7444
rect 6500 7108 6564 7172
rect 6684 7168 6748 7172
rect 6684 7112 6734 7168
rect 6734 7112 6748 7168
rect 6684 7108 6748 7112
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 5396 6972 5460 7036
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 5764 6896 5828 6900
rect 5764 6840 5778 6896
rect 5778 6840 5828 6896
rect 5764 6836 5828 6840
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 17612 6556 17676 6560
rect 17612 6500 17616 6556
rect 17616 6500 17672 6556
rect 17672 6500 17676 6556
rect 17612 6496 17676 6500
rect 17692 6556 17756 6560
rect 17692 6500 17696 6556
rect 17696 6500 17752 6556
rect 17752 6500 17756 6556
rect 17692 6496 17756 6500
rect 17772 6556 17836 6560
rect 17772 6500 17776 6556
rect 17776 6500 17832 6556
rect 17832 6500 17836 6556
rect 17772 6496 17836 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 8892 5748 8956 5812
rect 14964 5612 15028 5676
rect 3188 5476 3252 5540
rect 6684 5476 6748 5540
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 17612 5468 17676 5472
rect 17612 5412 17616 5468
rect 17616 5412 17672 5468
rect 17672 5412 17676 5468
rect 17612 5408 17676 5412
rect 17692 5468 17756 5472
rect 17692 5412 17696 5468
rect 17696 5412 17752 5468
rect 17752 5412 17756 5468
rect 17692 5408 17756 5412
rect 17772 5468 17836 5472
rect 17772 5412 17776 5468
rect 17776 5412 17832 5468
rect 17832 5412 17836 5468
rect 17772 5408 17836 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 5212 4856 5276 4860
rect 5212 4800 5262 4856
rect 5262 4800 5276 4856
rect 5212 4796 5276 4800
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 17612 4380 17676 4384
rect 17612 4324 17616 4380
rect 17616 4324 17672 4380
rect 17672 4324 17676 4380
rect 17612 4320 17676 4324
rect 17692 4380 17756 4384
rect 17692 4324 17696 4380
rect 17696 4324 17752 4380
rect 17752 4324 17756 4380
rect 17692 4320 17756 4324
rect 17772 4380 17836 4384
rect 17772 4324 17776 4380
rect 17776 4324 17832 4380
rect 17832 4324 17836 4380
rect 17772 4320 17836 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 11100 3768 11164 3772
rect 11100 3712 11150 3768
rect 11150 3712 11164 3768
rect 11100 3708 11164 3712
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 17612 3292 17676 3296
rect 17612 3236 17616 3292
rect 17616 3236 17672 3292
rect 17672 3236 17676 3292
rect 17612 3232 17676 3236
rect 17692 3292 17756 3296
rect 17692 3236 17696 3292
rect 17696 3236 17752 3292
rect 17752 3236 17756 3292
rect 17692 3232 17756 3236
rect 17772 3292 17836 3296
rect 17772 3236 17776 3292
rect 17776 3236 17832 3292
rect 17832 3236 17836 3292
rect 17772 3232 17836 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 9444 3028 9508 3092
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 15700 2484 15764 2548
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 17612 2204 17676 2208
rect 17612 2148 17616 2204
rect 17616 2148 17672 2204
rect 17672 2148 17676 2204
rect 17612 2144 17676 2148
rect 17692 2204 17756 2208
rect 17692 2148 17696 2204
rect 17696 2148 17752 2204
rect 17752 2148 17756 2204
rect 17692 2144 17756 2148
rect 17772 2204 17836 2208
rect 17772 2148 17776 2204
rect 17776 2148 17832 2204
rect 17832 2148 17836 2204
rect 17772 2144 17836 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
<< metal4 >>
rect 1944 16896 2264 17456
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 17440 2924 17456
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2604 16352 2924 17376
rect 6944 16896 7264 17456
rect 6944 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7264 16896
rect 5763 16556 5829 16557
rect 5763 16492 5764 16556
rect 5828 16492 5829 16556
rect 5763 16491 5829 16492
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 5395 15332 5461 15333
rect 5395 15268 5396 15332
rect 5460 15268 5461 15332
rect 5395 15267 5461 15268
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 5211 14924 5277 14925
rect 5211 14860 5212 14924
rect 5276 14860 5277 14924
rect 5211 14859 5277 14860
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 4107 13836 4173 13837
rect 4107 13772 4108 13836
rect 4172 13772 4173 13836
rect 4107 13771 4173 13772
rect 2604 13088 2924 13718
rect 3187 13292 3253 13293
rect 3187 13228 3188 13292
rect 3252 13228 3253 13292
rect 3187 13227 3253 13228
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 3190 5541 3250 13227
rect 4110 7445 4170 13771
rect 5027 12884 5093 12885
rect 5027 12820 5028 12884
rect 5092 12820 5093 12884
rect 5027 12819 5093 12820
rect 5030 9621 5090 12819
rect 5027 9620 5093 9621
rect 5027 9556 5028 9620
rect 5092 9556 5093 9620
rect 5027 9555 5093 9556
rect 4107 7444 4173 7445
rect 4107 7380 4108 7444
rect 4172 7380 4173 7444
rect 4107 7379 4173 7380
rect 3187 5540 3253 5541
rect 3187 5476 3188 5540
rect 3252 5476 3253 5540
rect 3187 5475 3253 5476
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 5214 4861 5274 14859
rect 5398 7037 5458 15267
rect 5395 7036 5461 7037
rect 5395 6972 5396 7036
rect 5460 6972 5461 7036
rect 5395 6971 5461 6972
rect 5766 6901 5826 16491
rect 6944 15808 7264 16832
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6944 14720 7264 15744
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 6944 13632 7264 14656
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 6944 12544 7264 13058
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 7604 17440 7924 17456
rect 7604 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7924 17440
rect 7604 16352 7924 17376
rect 11944 16896 12264 17456
rect 11944 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12264 16896
rect 8155 16692 8221 16693
rect 8155 16628 8156 16692
rect 8220 16628 8221 16692
rect 8155 16627 8221 16628
rect 7604 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7924 16352
rect 7604 15264 7924 16288
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7604 14176 7924 15200
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 7604 13088 7924 13718
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7604 12000 7924 13024
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7419 11932 7485 11933
rect 7419 11868 7420 11932
rect 7484 11868 7485 11932
rect 7419 11867 7485 11868
rect 7422 11525 7482 11867
rect 7419 11524 7485 11525
rect 7419 11460 7420 11524
rect 7484 11460 7485 11524
rect 7419 11459 7485 11460
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 6683 10980 6749 10981
rect 6683 10916 6684 10980
rect 6748 10916 6749 10980
rect 6683 10915 6749 10916
rect 6499 7852 6565 7853
rect 6499 7788 6500 7852
rect 6564 7788 6565 7852
rect 6499 7787 6565 7788
rect 6502 7173 6562 7787
rect 6686 7173 6746 10915
rect 6944 10368 7264 11392
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6944 9280 7264 10304
rect 7604 10912 7924 11936
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7604 9824 7924 10848
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7419 9756 7485 9757
rect 7419 9692 7420 9756
rect 7484 9692 7485 9756
rect 7419 9691 7485 9692
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 7422 9213 7482 9691
rect 7419 9212 7485 9213
rect 7419 9148 7420 9212
rect 7484 9148 7485 9212
rect 7419 9147 7485 9148
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6499 7172 6565 7173
rect 6499 7108 6500 7172
rect 6564 7108 6565 7172
rect 6499 7107 6565 7108
rect 6683 7172 6749 7173
rect 6683 7108 6684 7172
rect 6748 7108 6749 7172
rect 6683 7107 6749 7108
rect 5763 6900 5829 6901
rect 5763 6836 5764 6900
rect 5828 6836 5829 6900
rect 5763 6835 5829 6836
rect 6686 5541 6746 7107
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6683 5540 6749 5541
rect 6683 5476 6684 5540
rect 6748 5476 6749 5540
rect 6683 5475 6749 5476
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 5211 4860 5277 4861
rect 5211 4796 5212 4860
rect 5276 4796 5277 4860
rect 5211 4795 5277 4796
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 8954 7924 9760
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7604 7648 7924 8672
rect 8158 8669 8218 16627
rect 11944 15808 12264 16832
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 9627 15332 9693 15333
rect 9627 15268 9628 15332
rect 9692 15268 9693 15332
rect 9627 15267 9693 15268
rect 8891 13836 8957 13837
rect 8891 13772 8892 13836
rect 8956 13772 8957 13836
rect 8891 13771 8957 13772
rect 8339 12476 8405 12477
rect 8339 12412 8340 12476
rect 8404 12412 8405 12476
rect 8339 12411 8405 12412
rect 8342 9893 8402 12411
rect 8339 9892 8405 9893
rect 8339 9828 8340 9892
rect 8404 9828 8405 9892
rect 8339 9827 8405 9828
rect 8155 8668 8221 8669
rect 8155 8604 8156 8668
rect 8220 8604 8221 8668
rect 8155 8603 8221 8604
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 8894 5813 8954 13771
rect 9443 11116 9509 11117
rect 9443 11052 9444 11116
rect 9508 11052 9509 11116
rect 9443 11051 9509 11052
rect 8891 5812 8957 5813
rect 8891 5748 8892 5812
rect 8956 5748 8957 5812
rect 8891 5747 8957 5748
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 9446 3093 9506 11051
rect 9630 10709 9690 15267
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11944 13632 12264 14656
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 9811 11524 9877 11525
rect 9811 11460 9812 11524
rect 9876 11460 9877 11524
rect 9811 11459 9877 11460
rect 9627 10708 9693 10709
rect 9627 10644 9628 10708
rect 9692 10644 9693 10708
rect 9627 10643 9693 10644
rect 9814 8397 9874 11459
rect 11944 11456 12264 12480
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 10179 11388 10245 11389
rect 10179 11324 10180 11388
rect 10244 11324 10245 11388
rect 10179 11323 10245 11324
rect 10182 10981 10242 11323
rect 10179 10980 10245 10981
rect 10179 10916 10180 10980
rect 10244 10916 10245 10980
rect 10179 10915 10245 10916
rect 11099 10572 11165 10573
rect 11099 10508 11100 10572
rect 11164 10508 11165 10572
rect 11099 10507 11165 10508
rect 9811 8396 9877 8397
rect 9811 8332 9812 8396
rect 9876 8332 9877 8396
rect 9811 8331 9877 8332
rect 11102 3773 11162 10507
rect 11944 10368 12264 11392
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 11944 4928 12264 5952
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11099 3772 11165 3773
rect 11099 3708 11100 3772
rect 11164 3708 11165 3772
rect 11099 3707 11165 3708
rect 11944 3294 12264 3776
rect 9443 3092 9509 3093
rect 9443 3028 9444 3092
rect 9508 3028 9509 3092
rect 9443 3027 9509 3028
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 11944 2128 12264 2688
rect 12604 17440 12924 17456
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 16944 16896 17264 17456
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 13859 15332 13925 15333
rect 13859 15268 13860 15332
rect 13924 15268 13925 15332
rect 13859 15267 13925 15268
rect 14963 15332 15029 15333
rect 14963 15268 14964 15332
rect 15028 15268 15029 15332
rect 14963 15267 15029 15268
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 12604 13088 12924 13718
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12604 8954 12924 9760
rect 13862 9077 13922 15267
rect 13859 9076 13925 9077
rect 13859 9012 13860 9076
rect 13924 9012 13925 9076
rect 13859 9011 13925 9012
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 14966 5677 15026 15267
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13294 17264 13568
rect 15699 13156 15765 13157
rect 15699 13092 15700 13156
rect 15764 13092 15765 13156
rect 15699 13091 15765 13092
rect 15147 9756 15213 9757
rect 15147 9692 15148 9756
rect 15212 9692 15213 9756
rect 15147 9691 15213 9692
rect 15150 7989 15210 9691
rect 15147 7988 15213 7989
rect 15147 7924 15148 7988
rect 15212 7924 15213 7988
rect 15147 7923 15213 7924
rect 14963 5676 15029 5677
rect 14963 5612 14964 5676
rect 15028 5612 15029 5676
rect 14963 5611 15029 5612
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 15702 2549 15762 13091
rect 16944 13058 16986 13294
rect 17222 13058 17264 13294
rect 16803 12748 16869 12749
rect 16803 12684 16804 12748
rect 16868 12684 16869 12748
rect 16803 12683 16869 12684
rect 16806 12341 16866 12683
rect 16944 12544 17264 13058
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16803 12340 16869 12341
rect 16803 12276 16804 12340
rect 16868 12276 16869 12340
rect 16803 12275 16869 12276
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8294 17264 9216
rect 16944 8192 16986 8294
rect 17222 8192 17264 8294
rect 16944 8128 16952 8192
rect 17256 8128 17264 8192
rect 16944 8058 16986 8128
rect 17222 8058 17264 8128
rect 16944 7104 17264 8058
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3294 17264 3776
rect 16944 3058 16986 3294
rect 17222 3058 17264 3294
rect 16944 2752 17264 3058
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 15699 2548 15765 2549
rect 15699 2484 15700 2548
rect 15764 2484 15765 2548
rect 15699 2483 15765 2484
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 16944 2128 17264 2688
rect 17604 17440 17924 17456
rect 17604 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17924 17440
rect 17604 16352 17924 17376
rect 17604 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17924 16352
rect 17604 15264 17924 16288
rect 17604 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17924 15264
rect 17604 14176 17924 15200
rect 17604 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17924 14176
rect 17604 13954 17924 14112
rect 17604 13718 17646 13954
rect 17882 13718 17924 13954
rect 17604 13088 17924 13718
rect 17604 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17924 13088
rect 17604 12000 17924 13024
rect 17604 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17924 12000
rect 17604 10912 17924 11936
rect 17604 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17924 10912
rect 17604 9824 17924 10848
rect 17604 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17924 9824
rect 17604 8954 17924 9760
rect 17604 8736 17646 8954
rect 17882 8736 17924 8954
rect 17604 8672 17612 8736
rect 17676 8672 17692 8718
rect 17756 8672 17772 8718
rect 17836 8672 17852 8718
rect 17916 8672 17924 8736
rect 17604 7648 17924 8672
rect 17604 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17924 7648
rect 17604 6560 17924 7584
rect 17604 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17924 6560
rect 17604 5472 17924 6496
rect 17604 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17924 5472
rect 17604 4384 17924 5408
rect 17604 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17924 4384
rect 17604 3954 17924 4320
rect 17604 3718 17646 3954
rect 17882 3718 17924 3954
rect 17604 3296 17924 3718
rect 17604 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17924 3296
rect 17604 2208 17924 3232
rect 17604 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17924 2208
rect 17604 2128 17924 2144
<< via4 >>
rect 1986 13058 2222 13294
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1986 3058 2222 3294
rect 2646 13718 2882 13954
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 6986 13058 7222 13294
rect 7646 13718 7882 13954
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 2646 3718 2882 3954
rect 6986 3058 7222 3294
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 7646 3718 7882 3954
rect 11986 13058 12222 13294
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 11986 3058 12222 3294
rect 12646 13718 12882 13954
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 12646 3718 12882 3954
rect 16986 13058 17222 13294
rect 16986 8192 17222 8294
rect 16986 8128 17016 8192
rect 17016 8128 17032 8192
rect 17032 8128 17096 8192
rect 17096 8128 17112 8192
rect 17112 8128 17176 8192
rect 17176 8128 17192 8192
rect 17192 8128 17222 8192
rect 16986 8058 17222 8128
rect 16986 3058 17222 3294
rect 17646 13718 17882 13954
rect 17646 8736 17882 8954
rect 17646 8718 17676 8736
rect 17676 8718 17692 8736
rect 17692 8718 17756 8736
rect 17756 8718 17772 8736
rect 17772 8718 17836 8736
rect 17836 8718 17852 8736
rect 17852 8718 17882 8736
rect 17646 3718 17882 3954
<< metal5 >>
rect 1056 13954 18908 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 17646 13954
rect 17882 13718 18908 13954
rect 1056 13676 18908 13718
rect 1056 13294 18908 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 16986 13294
rect 17222 13058 18908 13294
rect 1056 13016 18908 13058
rect 1056 8954 18908 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 17646 8954
rect 17882 8718 18908 8954
rect 1056 8676 18908 8718
rect 1056 8294 18908 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 16986 8294
rect 17222 8058 18908 8294
rect 1056 8016 18908 8058
rect 1056 3954 18908 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 17646 3954
rect 17882 3718 18908 3954
rect 1056 3676 18908 3718
rect 1056 3294 18908 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 16986 3294
rect 17222 3058 18908 3294
rect 1056 3016 18908 3058
use sky130_ef_sc_hd__decap_12  FILLER_0_1_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_9
timestamp 1633347170
transform 1 0 1932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 1932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1633347170
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1633347170
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1633347170
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_33
timestamp 1633347170
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1633347170
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_45
timestamp 1633347170
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 1633347170
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 6348 0 -1 3264
box -38 -48 498 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_62
timestamp 1633347170
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1633347170
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69
timestamp 1633347170
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_53
timestamp 1633347170
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_49
timestamp 1633347170
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1633347170
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1633347170
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1633347170
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_77
timestamp 1633347170
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1633347170
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_86
timestamp 1633347170
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_94
timestamp 1633347170
transform 1 0 9752 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1633347170
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_90
timestamp 1633347170
transform 1 0 9384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_74
timestamp 1633347170
transform 1 0 7912 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 9292 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__o21a_1  _146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 10488 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 11500 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_118
timestamp 1633347170
transform 1 0 11960 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_108
timestamp 1633347170
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1633347170
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1633347170
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1633347170
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1633347170
transform 1 0 13064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_128
timestamp 1633347170
transform 1 0 12880 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 1633347170
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp 1633347170
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_133
timestamp 1633347170
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_120
timestamp 1633347170
transform 1 0 12144 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_130
timestamp 1633347170
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1633347170
transform 1 0 14260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1633347170
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _184_
timestamp 1633347170
transform 1 0 16100 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_157 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 15548 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_161
timestamp 1633347170
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_149
timestamp 1633347170
transform 1 0 14812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _183_
timestamp 1633347170
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _162_
timestamp 1633347170
transform 1 0 14720 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_145
timestamp 1633347170
transform 1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1633347170
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1633347170
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_169
timestamp 1633347170
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1633347170
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1633347170
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 16928 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_184
timestamp 1633347170
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1633347170
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_179
timestamp 1633347170
transform 1 0 17572 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 1633347170
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_187
timestamp 1633347170
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1633347170
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1633347170
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1633347170
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_22
timestamp 1633347170
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_10
timestamp 1633347170
transform 1 0 2024 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1633347170
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 5428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3772 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_39
timestamp 1633347170
transform 1 0 4692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1633347170
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1633347170
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1633347170
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _290_
timestamp 1633347170
transform 1 0 8924 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1633347170
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1633347170
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1633347170
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a221oi_4  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 11040 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_141
timestamp 1633347170
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_129
timestamp 1633347170
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_137
timestamp 1633347170
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1633347170
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 14628 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 15456 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1633347170
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_180
timestamp 1633347170
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1633347170
transform 1 0 18032 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1633347170
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 1472 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _194_
timestamp 1633347170
transform 1 0 2116 0 -1 4352
box -38 -48 498 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_16
timestamp 1633347170
transform 1 0 2576 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1633347170
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1633347170
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 4048 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_28
timestamp 1633347170
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_57
timestamp 1633347170
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_71
timestamp 1633347170
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1633347170
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1633347170
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_65
timestamp 1633347170
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1633347170
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _161_
timestamp 1633347170
transform 1 0 8004 0 -1 4352
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_94
timestamp 1633347170
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_82
timestamp 1633347170
transform 1 0 8648 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _284_
timestamp 1633347170
transform 1 0 11500 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_106
timestamp 1633347170
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1633347170
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_133
timestamp 1633347170
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_145
timestamp 1633347170
transform 1 0 14444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_157
timestamp 1633347170
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_165
timestamp 1633347170
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _182_
timestamp 1633347170
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 18032 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_175
timestamp 1633347170
transform 1 0 17204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_183
timestamp 1633347170
transform 1 0 17940 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_179
timestamp 1633347170
transform 1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1633347170
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1633347170
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _292_
timestamp 1633347170
transform 1 0 1380 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1633347170
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _137_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3772 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_47
timestamp 1633347170
transform 1 0 5428 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_24
timestamp 1633347170
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1633347170
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 6992 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_8  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 5980 0 1 4352
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_71
timestamp 1633347170
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _225_
timestamp 1633347170
transform 1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_85
timestamp 1633347170
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_91
timestamp 1633347170
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1633347170
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1633347170
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _295_
timestamp 1633347170
transform 1 0 11592 0 1 4352
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_99
timestamp 1633347170
transform 1 0 10212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_111
timestamp 1633347170
transform 1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_134
timestamp 1633347170
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1633347170
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1633347170
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _300_
timestamp 1633347170
transform 1 0 15180 0 1 4352
box -38 -48 1970 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_174
timestamp 1633347170
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_186
timestamp 1633347170
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1633347170
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 1380 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _193_
timestamp 1633347170
transform 1 0 2208 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_19
timestamp 1633347170
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1633347170
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _280_
timestamp 1633347170
transform 1 0 3680 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_27
timestamp 1633347170
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 7268 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_65
timestamp 1633347170
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1633347170
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_48
timestamp 1633347170
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1633347170
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_86
timestamp 1633347170
transform 1 0 9016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_74
timestamp 1633347170
transform 1 0 7912 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _179_
timestamp 1633347170
transform 1 0 11500 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1633347170
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_98
timestamp 1633347170
transform 1 0 10120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1633347170
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1633347170
transform 1 0 12144 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_135
timestamp 1633347170
transform 1 0 13524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_123
timestamp 1633347170
transform 1 0 12420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 1633347170
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_147
timestamp 1633347170
transform 1 0 14628 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  fanout31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 15640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1633347170
transform 1 0 16008 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_155
timestamp 1633347170
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1633347170
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_189
timestamp 1633347170
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_181
timestamp 1633347170
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1633347170
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1633347170
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o21ba_1  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 2300 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3036 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1633347170
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1633347170
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1633347170
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_12
timestamp 1633347170
transform 1 0 2208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1633347170
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1633347170
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1633347170
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1633347170
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _172_
timestamp 1633347170
transform 1 0 3956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_27
timestamp 1633347170
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1633347170
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1633347170
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_34
timestamp 1633347170
transform 1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_46
timestamp 1633347170
transform 1 0 5336 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_34
timestamp 1633347170
transform 1 0 4232 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _282_
timestamp 1633347170
transform 1 0 5428 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _297_
timestamp 1633347170
transform 1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  _186_
timestamp 1633347170
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _176_
timestamp 1633347170
transform 1 0 7360 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_2  _294_
timestamp 1633347170
transform 1 0 7544 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_64
timestamp 1633347170
transform 1 0 6992 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_67
timestamp 1633347170
transform 1 0 7268 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1633347170
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__and4_2  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _188_
timestamp 1633347170
transform 1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_85
timestamp 1633347170
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_91
timestamp 1633347170
transform 1 0 9476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_91
timestamp 1633347170
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1633347170
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1633347170
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _222_
timestamp 1633347170
transform 1 0 11776 0 1 5440
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1633347170
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_99
timestamp 1633347170
transform 1 0 10212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1633347170
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_115
timestamp 1633347170
transform 1 0 11684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_103
timestamp 1633347170
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_111
timestamp 1633347170
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1633347170
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _207_
timestamp 1633347170
transform 1 0 13708 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_141
timestamp 1633347170
transform 1 0 14076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1633347170
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1633347170
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_123
timestamp 1633347170
transform 1 0 12420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1633347170
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_135
timestamp 1633347170
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1633347170
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_153
timestamp 1633347170
transform 1 0 15180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_159
timestamp 1633347170
transform 1 0 15732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _166_
timestamp 1633347170
transform 1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1633347170
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_153
timestamp 1633347170
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1633347170
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1633347170
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1633347170
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1633347170
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_181
timestamp 1633347170
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_189
timestamp 1633347170
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_185
timestamp 1633347170
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_183
timestamp 1633347170
transform 1 0 17940 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_171
timestamp 1633347170
transform 1 0 16836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1633347170
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1633347170
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1633347170
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1633347170
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1633347170
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1633347170
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1633347170
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1633347170
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1633347170
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1633347170
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1633347170
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1633347170
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1633347170
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1633347170
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1633347170
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1633347170
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1633347170
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1633347170
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1633347170
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1633347170
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1633347170
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1633347170
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_165
timestamp 1633347170
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1633347170
transform 1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1633347170
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_186
timestamp 1633347170
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_179
timestamp 1633347170
transform 1 0 17572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1633347170
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_173
timestamp 1633347170
transform 1 0 17020 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1633347170
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1633347170
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1633347170
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _175_
timestamp 1633347170
transform 1 0 5244 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_39
timestamp 1633347170
transform 1 0 4692 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1633347170
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _228_
timestamp 1633347170
transform 1 0 6348 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_64
timestamp 1633347170
transform 1 0 6992 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_70
timestamp 1633347170
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1633347170
transform 1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1633347170
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_87
timestamp 1633347170
transform 1 0 9108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_75
timestamp 1633347170
transform 1 0 8004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _141_
timestamp 1633347170
transform 1 0 11960 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_99
timestamp 1633347170
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_117
timestamp 1633347170
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1633347170
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 1633347170
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1633347170
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_136
timestamp 1633347170
transform 1 0 13616 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_124
timestamp 1633347170
transform 1 0 12512 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_148
timestamp 1633347170
transform 1 0 14720 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_160
timestamp 1633347170
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1633347170
transform 1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1633347170
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_189
timestamp 1633347170
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_181
timestamp 1633347170
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_185
timestamp 1633347170
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1633347170
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1633347170
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1633347170
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_21
timestamp 1633347170
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1633347170
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1633347170
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_15
timestamp 1633347170
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1633347170
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1633347170
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1633347170
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1633347170
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _234_
timestamp 1633347170
transform 1 0 6256 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_62
timestamp 1633347170
transform 1 0 6808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_53
timestamp 1633347170
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _171_
timestamp 1633347170
transform 1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1633347170
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_93
timestamp 1633347170
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1633347170
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_74
timestamp 1633347170
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1633347170
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1633347170
transform 1 0 10948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_100
timestamp 1633347170
transform 1 0 10304 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_110
timestamp 1633347170
transform 1 0 11224 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_106
timestamp 1633347170
transform 1 0 10856 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp 1633347170
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1633347170
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_122
timestamp 1633347170
transform 1 0 12328 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1633347170
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1633347170
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1633347170
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1633347170
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_189
timestamp 1633347170
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1633347170
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_23
timestamp 1633347170
transform 1 0 3220 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1633347170
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_15
timestamp 1633347170
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1633347170
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3404 0 -1 8704
box -38 -48 498 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_42
timestamp 1633347170
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1633347170
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_1  _150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 6348 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1633347170
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1633347170
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_90
timestamp 1633347170
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_78
timestamp 1633347170
transform 1 0 8280 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1633347170
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1633347170
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1633347170
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1633347170
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1633347170
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _229_
timestamp 1633347170
transform 1 0 13708 0 -1 8704
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1633347170
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_156
timestamp 1633347170
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_144
timestamp 1633347170
transform 1 0 14352 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _165_
timestamp 1633347170
transform 1 0 17664 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1633347170
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_186
timestamp 1633347170
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1633347170
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_177
timestamp 1633347170
transform 1 0 17388 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1633347170
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1633347170
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1633347170
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1633347170
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1633347170
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1633347170
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1633347170
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1633347170
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1633347170
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _142_
timestamp 1633347170
transform 1 0 7636 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 6256 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_64
timestamp 1633347170
transform 1 0 6992 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_70
timestamp 1633347170
transform 1 0 7544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_53
timestamp 1633347170
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _174_
timestamp 1633347170
transform 1 0 8924 0 1 8704
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_92
timestamp 1633347170
transform 1 0 9568 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1633347170
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1633347170
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_104
timestamp 1633347170
transform 1 0 10672 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_116
timestamp 1633347170
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _286_
timestamp 1633347170
transform 1 0 12144 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_141
timestamp 1633347170
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1633347170
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  _248_
timestamp 1633347170
transform 1 0 14904 0 1 8704
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_161
timestamp 1633347170
transform 1 0 15916 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_149
timestamp 1633347170
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_173
timestamp 1633347170
transform 1 0 17020 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_189
timestamp 1633347170
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_185
timestamp 1633347170
transform 1 0 18124 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1633347170
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1633347170
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1633347170
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1633347170
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_21
timestamp 1633347170
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_9
timestamp 1633347170
transform 1 0 1932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1633347170
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1633347170
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_3
timestamp 1633347170
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _221_
timestamp 1633347170
transform 1 0 4324 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _274_
timestamp 1633347170
transform 1 0 4968 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_29
timestamp 1633347170
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_41
timestamp 1633347170
transform 1 0 4876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1633347170
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_33
timestamp 1633347170
transform 1 0 4140 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _148_
timestamp 1633347170
transform 1 0 5060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1633347170
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _195_
timestamp 1633347170
transform 1 0 7176 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_2  _301_
timestamp 1633347170
transform 1 0 6440 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_49
timestamp 1633347170
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1633347170
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1633347170
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_62
timestamp 1633347170
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1633347170
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _296_
timestamp 1633347170
transform 1 0 8556 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_79
timestamp 1633347170
transform 1 0 8372 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1633347170
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_73
timestamp 1633347170
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1633347170
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1633347170
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _279_
timestamp 1633347170
transform 1 0 10580 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_97
timestamp 1633347170
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1633347170
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1633347170
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp 1633347170
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1633347170
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_124
timestamp 1633347170
transform 1 0 12512 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1633347170
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1633347170
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _214_
timestamp 1633347170
transform 1 0 13432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_138
timestamp 1633347170
transform 1 0 13800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_135
timestamp 1633347170
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_142
timestamp 1633347170
transform 1 0 14168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1633347170
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_132
timestamp 1633347170
transform 1 0 13248 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_1  _212_
timestamp 1633347170
transform 1 0 14260 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_123
timestamp 1633347170
transform 1 0 12420 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1633347170
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _215_
timestamp 1633347170
transform 1 0 15640 0 1 9792
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_147
timestamp 1633347170
transform 1 0 14628 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1633347170
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_165
timestamp 1633347170
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_159
timestamp 1633347170
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1633347170
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1633347170
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1633347170
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__and4_2  _155_
timestamp 1633347170
transform 1 0 17020 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_181
timestamp 1633347170
transform 1 0 17756 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1633347170
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1633347170
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 1633347170
transform 1 0 18032 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_181
timestamp 1633347170
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_189
timestamp 1633347170
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1633347170
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1633347170
transform 1 0 2668 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_20
timestamp 1633347170
transform 1 0 2944 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_15
timestamp 1633347170
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1633347170
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1633347170
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1633347170
transform 1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_42
timestamp 1633347170
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_30
timestamp 1633347170
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_26
timestamp 1633347170
transform 1 0 3496 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1633347170
transform 1 0 7452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1633347170
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1633347170
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1633347170
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_84
timestamp 1633347170
transform 1 0 8832 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_72
timestamp 1633347170
transform 1 0 7728 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1633347170
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_96
timestamp 1633347170
transform 1 0 9936 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 1633347170
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1633347170
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1633347170
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1633347170
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _177_
timestamp 1633347170
transform 1 0 14904 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_156
timestamp 1633347170
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_149
timestamp 1633347170
transform 1 0 14812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _200_
timestamp 1633347170
transform 1 0 17940 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _218_
timestamp 1633347170
transform 1 0 17204 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_169
timestamp 1633347170
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_188
timestamp 1633347170
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_181
timestamp 1633347170
transform 1 0 17756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1633347170
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1633347170
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1633347170
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1633347170
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1633347170
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _235_
timestamp 1633347170
transform 1 0 4508 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_44
timestamp 1633347170
transform 1 0 5152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1633347170
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1633347170
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_68
timestamp 1633347170
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_56
timestamp 1633347170
transform 1 0 6256 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _190_
timestamp 1633347170
transform 1 0 9568 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _181_
timestamp 1633347170
transform 1 0 8924 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 1633347170
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1633347170
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _288_
timestamp 1633347170
transform 1 0 10304 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_98
timestamp 1633347170
transform 1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _277_
timestamp 1633347170
transform 1 0 14076 0 1 10880
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_123
timestamp 1633347170
transform 1 0 12420 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1633347170
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_135
timestamp 1633347170
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1633347170
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_161
timestamp 1633347170
transform 1 0 15916 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _153_
timestamp 1633347170
transform 1 0 18124 0 1 10880
box -38 -48 498 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_173
timestamp 1633347170
transform 1 0 17020 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1633347170
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_4  _152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 1840 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_7
timestamp 1633347170
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_3
timestamp 1633347170
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1633347170
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_38
timestamp 1633347170
transform 1 0 4600 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_26
timestamp 1633347170
transform 1 0 3496 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_1  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 6992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _219_
timestamp 1633347170
transform 1 0 6348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_50
timestamp 1633347170
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_70
timestamp 1633347170
transform 1 0 7544 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1633347170
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_82
timestamp 1633347170
transform 1 0 8648 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_94
timestamp 1633347170
transform 1 0 9752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _231_
timestamp 1633347170
transform 1 0 10212 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_106
timestamp 1633347170
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_98
timestamp 1633347170
transform 1 0 10120 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_113
timestamp 1633347170
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1633347170
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _299_
timestamp 1633347170
transform 1 0 12236 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1633347170
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1633347170
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_146
timestamp 1633347170
transform 1 0 14536 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_158
timestamp 1633347170
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1633347170
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_189
timestamp 1633347170
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1633347170
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1633347170
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1633347170
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _230_
timestamp 1633347170
transform 1 0 2024 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _233_
timestamp 1633347170
transform 1 0 2944 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1633347170
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_9
timestamp 1633347170
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_16
timestamp 1633347170
transform 1 0 2576 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1633347170
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1633347170
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1633347170
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1633347170
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1633347170
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _164_
timestamp 1633347170
transform 1 0 6072 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1633347170
transform 1 0 7268 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_61
timestamp 1633347170
transform 1 0 6716 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_70
timestamp 1633347170
transform 1 0 7544 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_53
timestamp 1633347170
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _158_
timestamp 1633347170
transform 1 0 9568 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _232_
timestamp 1633347170
transform 1 0 8924 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1633347170
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1633347170
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 10304 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_108
timestamp 1633347170
transform 1 0 11040 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_97
timestamp 1633347170
transform 1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _154_
timestamp 1633347170
transform 1 0 14076 0 1 11968
box -38 -48 498 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_120
timestamp 1633347170
transform 1 0 12144 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_132
timestamp 1633347170
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1633347170
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_158
timestamp 1633347170
transform 1 0 15640 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_146
timestamp 1633347170
transform 1 0 14536 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_170
timestamp 1633347170
transform 1 0 16744 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_182
timestamp 1633347170
transform 1 0 17848 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1633347170
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _276_
timestamp 1633347170
transform 1 0 2576 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_14
timestamp 1633347170
transform 1 0 2392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1633347170
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_6
timestamp 1633347170
transform 1 0 1656 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_23
timestamp 1633347170
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1633347170
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1633347170
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1633347170
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1633347170
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_44
timestamp 1633347170
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_32
timestamp 1633347170
transform 1 0 4048 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_36
timestamp 1633347170
transform 1 0 4416 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1633347170
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1633347170
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _180_
timestamp 1633347170
transform 1 0 6992 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1633347170
transform 1 0 6256 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _283_
timestamp 1633347170
transform 1 0 7636 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 1633347170
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_71
timestamp 1633347170
transform 1 0 7636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_59
timestamp 1633347170
transform 1 0 6532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_63
timestamp 1633347170
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_48
timestamp 1633347170
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1633347170
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1633347170
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_91
timestamp 1633347170
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1633347170
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1633347170
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1633347170
transform 1 0 10580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_97
timestamp 1633347170
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_118
timestamp 1633347170
transform 1 0 11960 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_106
timestamp 1633347170
transform 1 0 10856 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1633347170
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1633347170
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_103
timestamp 1633347170
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1633347170
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _198_
timestamp 1633347170
transform 1 0 14076 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1633347170
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_130
timestamp 1633347170
transform 1 0 13064 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1633347170
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_136
timestamp 1633347170
transform 1 0 13616 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_137
timestamp 1633347170
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1633347170
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _293_
timestamp 1633347170
transform 1 0 15548 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _281_
timestamp 1633347170
transform 1 0 14720 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  _140_
timestamp 1633347170
transform 1 0 14996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_148
timestamp 1633347170
transform 1 0 14720 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_145
timestamp 1633347170
transform 1 0 14444 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_178
timestamp 1633347170
transform 1 0 17480 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1633347170
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1633347170
transform 1 0 18032 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1633347170
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1633347170
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_181
timestamp 1633347170
transform 1 0 17756 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1633347170
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _291_
timestamp 1633347170
transform 1 0 2484 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1633347170
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_13
timestamp 1633347170
transform 1 0 2300 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 1633347170
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1633347170
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1633347170
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1633347170
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _278_
timestamp 1633347170
transform 1 0 7176 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_61
timestamp 1633347170
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1633347170
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1633347170
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1633347170
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _227_
timestamp 1633347170
transform 1 0 6808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1633347170
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_86
timestamp 1633347170
transform 1 0 9016 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1633347170
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1633347170
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_98
timestamp 1633347170
transform 1 0 10120 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1633347170
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _287_
timestamp 1633347170
transform 1 0 13800 0 -1 14144
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1633347170
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_137
timestamp 1633347170
transform 1 0 13708 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1633347170
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_158
timestamp 1633347170
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1633347170
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 1633347170
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_181
timestamp 1633347170
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1633347170
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1633347170
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _226_
timestamp 1633347170
transform 1 0 2760 0 1 14144
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1633347170
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1633347170
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_15
timestamp 1633347170
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1633347170
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1633347170
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_25
timestamp 1633347170
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1633347170
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1633347170
transform 1 0 6164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1633347170
transform 1 0 6440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_53
timestamp 1633347170
transform 1 0 5980 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_61
timestamp 1633347170
transform 1 0 6716 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1633347170
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_73
timestamp 1633347170
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1633347170
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1633347170
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _213_
timestamp 1633347170
transform 1 0 12052 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1633347170
transform 1 0 11776 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_109
timestamp 1633347170
transform 1 0 11132 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1633347170
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_115
timestamp 1633347170
transform 1 0 11684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_132
timestamp 1633347170
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1633347170
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_124
timestamp 1633347170
transform 1 0 12512 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _191_
timestamp 1633347170
transform 1 0 13432 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1633347170
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1633347170
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1633347170
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_165
timestamp 1633347170
transform 1 0 16284 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 17020 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1633347170
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_189
timestamp 1633347170
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1633347170
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1633347170
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1633347170
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1633347170
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1633347170
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1633347170
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1633347170
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1633347170
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1633347170
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1633347170
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1633347170
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1633347170
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1633347170
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _159_
timestamp 1633347170
transform 1 0 11592 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1633347170
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_113
timestamp 1633347170
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_105
timestamp 1633347170
transform 1 0 10764 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1633347170
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _273_
timestamp 1633347170
transform 1 0 12328 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_121
timestamp 1633347170
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_142
timestamp 1633347170
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1633347170
transform 1 0 15180 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_156
timestamp 1633347170
transform 1 0 15456 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_146
timestamp 1633347170
transform 1 0 14536 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _163_
timestamp 1633347170
transform 1 0 14628 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _138_
timestamp 1633347170
transform 1 0 17664 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1633347170
transform 1 0 17296 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_183
timestamp 1633347170
transform 1 0 17940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_169
timestamp 1633347170
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_178
timestamp 1633347170
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_189
timestamp 1633347170
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_175
timestamp 1633347170
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1633347170
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1633347170
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_21
timestamp 1633347170
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_9
timestamp 1633347170
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1633347170
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1633347170
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _167_
timestamp 1633347170
transform 1 0 4784 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _259_
timestamp 1633347170
transform 1 0 3772 0 1 15232
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_45
timestamp 1633347170
transform 1 0 5244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1633347170
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1633347170
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_69
timestamp 1633347170
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_57
timestamp 1633347170
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1633347170
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1633347170
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1633347170
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _302_
timestamp 1633347170
transform 1 0 10672 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_97
timestamp 1633347170
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_103
timestamp 1633347170
transform 1 0 10580 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _224_
timestamp 1633347170
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _285_
timestamp 1633347170
transform 1 0 14076 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_132
timestamp 1633347170
transform 1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_124
timestamp 1633347170
transform 1 0 12512 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1633347170
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_161
timestamp 1633347170
transform 1 0 15916 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_173
timestamp 1633347170
transform 1 0 17020 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_189
timestamp 1633347170
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_185
timestamp 1633347170
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1633347170
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _187_
timestamp 1633347170
transform 1 0 2944 0 -1 16320
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1633347170
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_19
timestamp 1633347170
transform 1 0 2852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_15
timestamp 1633347170
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1633347170
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1633347170
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1633347170
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1633347170
transform 1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1633347170
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1633347170
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1633347170
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1633347170
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _275_
timestamp 1633347170
transform 1 0 7728 0 -1 16320
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_92
timestamp 1633347170
transform 1 0 9568 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 1633347170
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_104
timestamp 1633347170
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1633347170
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_1  _189_
timestamp 1633347170
transform 1 0 12420 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _272_
timestamp 1633347170
transform 1 0 13156 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_121
timestamp 1633347170
transform 1 0 12236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _211_
timestamp 1633347170
transform 1 0 14996 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1633347170
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1633347170
transform 1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_162
timestamp 1633347170
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_154
timestamp 1633347170
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__xor2_1  _169_
timestamp 1633347170
transform 1 0 16652 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_184
timestamp 1633347170
transform 1 0 18032 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_176
timestamp 1633347170
transform 1 0 17296 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1633347170
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1633347170
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1633347170
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_12
timestamp 1633347170
transform 1 0 2208 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1633347170
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1633347170
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1633347170
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1633347170
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1633347170
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1633347170
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1633347170
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1633347170
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1633347170
transform 1 0 3956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_29
timestamp 1633347170
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_24
timestamp 1633347170
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1633347170
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_29
timestamp 1633347170
transform 1 0 3772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_2  _145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633347170
transform 1 0 4140 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1633347170
transform 1 0 4508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _160_
timestamp 1633347170
transform 1 0 4784 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_40
timestamp 1633347170
transform 1 0 4784 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_57
timestamp 1633347170
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_65
timestamp 1633347170
transform 1 0 7084 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_64
timestamp 1633347170
transform 1 0 6992 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_52
timestamp 1633347170
transform 1 0 5888 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_48
timestamp 1633347170
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1633347170
transform 1 0 6532 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1633347170
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_77
timestamp 1633347170
transform 1 0 8188 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1633347170
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_93
timestamp 1633347170
transform 1 0 9660 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_83
timestamp 1633347170
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_85
timestamp 1633347170
transform 1 0 8924 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_76
timestamp 1633347170
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1633347170
transform 1 0 9752 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1633347170
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1633347170
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1633347170
transform 1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1633347170
transform 1 0 10028 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_112
timestamp 1633347170
transform 1 0 11408 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_100
timestamp 1633347170
transform 1 0 10304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_113
timestamp 1633347170
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_101
timestamp 1633347170
transform 1 0 10396 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1633347170
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1633347170
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_124
timestamp 1633347170
transform 1 0 12512 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1633347170
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_130
timestamp 1633347170
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_121
timestamp 1633347170
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1633347170
transform 1 0 12788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1633347170
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1633347170
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1633347170
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_138
timestamp 1633347170
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__and2_1  _173_
timestamp 1633347170
transform 1 0 14076 0 1 16320
box -38 -48 498 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_126
timestamp 1633347170
transform 1 0 12696 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_141
timestamp 1633347170
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_158
timestamp 1633347170
transform 1 0 15640 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_146
timestamp 1633347170
transform 1 0 14536 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_163
timestamp 1633347170
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_153
timestamp 1633347170
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1633347170
transform 1 0 15548 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1633347170
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_175
timestamp 1633347170
transform 1 0 17204 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 1633347170
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1633347170
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _185_
timestamp 1633347170
transform 1 0 16744 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_177
timestamp 1633347170
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1633347170
transform 1 0 18032 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1633347170
transform 1 0 17664 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_183
timestamp 1633347170
transform 1 0 17940 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1633347170
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1633347170
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_186
timestamp 1633347170
transform 1 0 18216 0 -1 17408
box -38 -48 406 592
<< labels >>
flabel metal4 s 2604 2128 2924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7604 2128 7924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12604 2128 12924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17604 2128 17924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3676 18908 3996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8676 18908 8996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 13676 18908 13996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6944 2128 7264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11944 2128 12264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 16944 2128 17264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3016 18908 3336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8016 18908 8336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 13016 18908 13336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 19200 8 20000 128 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 19200 6128 20000 6248 0 FreeSans 480 0 0 0 count[0]
port 3 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 count[10]
port 4 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 count[11]
port 5 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 count[12]
port 6 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 count[13]
port 7 nsew signal tristate
flabel metal2 s 18050 19200 18106 20000 0 FreeSans 224 90 0 0 count[14]
port 8 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 count[15]
port 9 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 count[1]
port 10 nsew signal tristate
flabel metal2 s 15474 19200 15530 20000 0 FreeSans 224 90 0 0 count[2]
port 11 nsew signal tristate
flabel metal3 s 19200 18368 20000 18488 0 FreeSans 480 0 0 0 count[3]
port 12 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 count[4]
port 13 nsew signal tristate
flabel metal2 s 3882 19200 3938 20000 0 FreeSans 224 90 0 0 count[5]
port 14 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 count[6]
port 15 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 count[7]
port 16 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 count[8]
port 17 nsew signal tristate
flabel metal2 s 6458 19200 6514 20000 0 FreeSans 224 90 0 0 count[9]
port 18 nsew signal tristate
flabel metal3 s 19200 3408 20000 3528 0 FreeSans 480 0 0 0 enable
port 19 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 inputData[0]
port 20 nsew signal input
flabel metal3 s 19200 12248 20000 12368 0 FreeSans 480 0 0 0 inputData[1]
port 21 nsew signal input
flabel metal3 s 19200 15648 20000 15768 0 FreeSans 480 0 0 0 inputData[2]
port 22 nsew signal input
flabel metal2 s 9678 19200 9734 20000 0 FreeSans 224 90 0 0 inputData[3]
port 23 nsew signal input
flabel metal2 s 12254 19200 12310 20000 0 FreeSans 224 90 0 0 inputData[4]
port 24 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 inputData[5]
port 25 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 inputData[6]
port 26 nsew signal input
flabel metal2 s 662 19200 718 20000 0 FreeSans 224 90 0 0 inputData[7]
port 27 nsew signal input
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 reset
port 28 nsew signal input
rlabel metal1 9982 17408 9982 17408 0 VGND
rlabel metal1 9982 16864 9982 16864 0 VPWR
rlabel via3 16859 12716 16859 12716 0 _000_
rlabel metal2 6578 14824 6578 14824 0 _001_
rlabel metal1 5152 13838 5152 13838 0 _002_
rlabel metal1 13294 3162 13294 3162 0 _003_
rlabel metal1 4837 12886 4837 12886 0 _004_
rlabel metal1 10212 16422 10212 16422 0 _005_
rlabel metal1 2254 6154 2254 6154 0 _006_
rlabel metal2 9798 8942 9798 8942 0 _007_
rlabel metal1 8050 8602 8050 8602 0 _008_
rlabel metal2 10718 13022 10718 13022 0 _009_
rlabel metal2 15318 14297 15318 14297 0 _010_
rlabel metal1 4232 10710 4232 10710 0 _011_
rlabel metal1 13163 4182 13163 4182 0 _012_
rlabel metal1 13938 15368 13938 15368 0 _013_
rlabel metal1 12052 13430 12052 13430 0 _014_
rlabel metal2 15226 13163 15226 13163 0 _015_
rlabel metal2 1794 10421 1794 10421 0 _016_
rlabel metal1 11047 2346 11047 2346 0 _017_
rlabel metal2 13754 5916 13754 5916 0 _018_
rlabel metal1 16928 6834 16928 6834 0 _019_
rlabel via2 13846 13243 13846 13243 0 _020_
rlabel via2 9154 2533 9154 2533 0 _021_
rlabel metal1 11960 5270 11960 5270 0 _022_
rlabel metal2 12466 9044 12466 9044 0 _023_
rlabel metal2 17526 3859 17526 3859 0 _024_
rlabel metal1 6401 6358 6401 6358 0 _025_
rlabel metal1 17165 3434 17165 3434 0 _026_
rlabel metal1 6578 17238 6578 17238 0 _027_
rlabel metal1 15686 15878 15686 15878 0 _028_
rlabel metal1 6663 9622 6663 9622 0 _029_
rlabel metal1 11362 15368 11362 15368 0 _030_
rlabel metal3 8418 14484 8418 14484 0 _031_
rlabel metal1 4048 16490 4048 16490 0 _032_
rlabel metal2 13018 13821 13018 13821 0 _033_
rlabel metal1 5796 8058 5796 8058 0 _034_
rlabel metal1 6072 15946 6072 15946 0 _035_
rlabel metal2 8970 12852 8970 12852 0 _036_
rlabel metal1 13386 11186 13386 11186 0 _037_
rlabel metal1 4048 12682 4048 12682 0 _038_
rlabel metal2 11178 9282 11178 9282 0 _039_
rlabel metal2 4002 6256 4002 6256 0 _040_
rlabel metal1 14858 12716 14858 12716 0 _041_
rlabel metal1 13340 15674 13340 15674 0 _042_
rlabel metal1 8556 12750 8556 12750 0 _043_
rlabel metal2 11822 3961 11822 3961 0 _044_
rlabel via2 14398 15419 14398 15419 0 _045_
rlabel metal2 11086 7803 11086 7803 0 _046_
rlabel metal1 14805 13702 14805 13702 0 _047_
rlabel metal1 3956 5882 3956 5882 0 _048_
rlabel metal1 9568 2346 9568 2346 0 _049_
rlabel metal1 10672 2890 10672 2890 0 _050_
rlabel via1 3542 13821 3542 13821 0 _051_
rlabel metal2 1702 4828 1702 4828 0 _052_
rlabel metal2 15870 13804 15870 13804 0 _053_
rlabel metal2 10166 6052 10166 6052 0 _054_
rlabel metal2 7498 5372 7498 5372 0 _055_
rlabel metal1 15180 2890 15180 2890 0 _056_
rlabel metal1 6164 12614 6164 12614 0 _057_
rlabel via2 15778 3451 15778 3451 0 _058_
rlabel metal2 13018 9384 13018 9384 0 _059_
rlabel metal2 13846 5423 13846 5423 0 _060_
rlabel metal1 17342 15878 17342 15878 0 _061_
rlabel metal1 11132 15402 11132 15402 0 _062_
rlabel metal1 8004 3978 8004 3978 0 _063_
rlabel metal2 1886 3264 1886 3264 0 _064_
rlabel metal1 17158 14858 17158 14858 0 _065_
rlabel metal1 2162 11764 2162 11764 0 _066_
rlabel metal2 7498 12478 7498 12478 0 _067_
rlabel metal1 15134 13430 15134 13430 0 _068_
rlabel metal1 7590 7514 7590 7514 0 _069_
rlabel metal1 2622 13260 2622 13260 0 _070_
rlabel metal2 2438 11900 2438 11900 0 _071_
rlabel metal2 2346 12478 2346 12478 0 _072_
rlabel metal2 13202 7004 13202 7004 0 _073_
rlabel metal1 11408 3162 11408 3162 0 _074_
rlabel metal2 1426 4233 1426 4233 0 _075_
rlabel metal2 1702 3570 1702 3570 0 _076_
rlabel metal1 2576 11730 2576 11730 0 _077_
rlabel metal2 3726 5457 3726 5457 0 _078_
rlabel metal1 1748 3706 1748 3706 0 _079_
rlabel metal2 14766 14790 14766 14790 0 _080_
rlabel metal1 16054 11322 16054 11322 0 _081_
rlabel metal1 11500 15130 11500 15130 0 _082_
rlabel metal1 12558 15980 12558 15980 0 _083_
rlabel metal2 15410 4947 15410 4947 0 _084_
rlabel metal2 9614 15300 9614 15300 0 _085_
rlabel metal1 5014 15572 5014 15572 0 _086_
rlabel metal1 5750 17170 5750 17170 0 _087_
rlabel metal3 6785 16660 6785 16660 0 _088_
rlabel metal1 18078 2958 18078 2958 0 _089_
rlabel metal1 18170 4046 18170 4046 0 _090_
rlabel metal2 15134 10047 15134 10047 0 _091_
rlabel metal1 16836 5678 16836 5678 0 _092_
rlabel metal2 16790 4131 16790 4131 0 _093_
rlabel metal1 17250 16014 17250 16014 0 _094_
rlabel metal1 16652 2958 16652 2958 0 _095_
rlabel metal2 8786 7412 8786 7412 0 _096_
rlabel metal1 11914 16762 11914 16762 0 _097_
rlabel metal1 12190 10574 12190 10574 0 _098_
rlabel metal2 15226 8432 15226 8432 0 _099_
rlabel metal4 15180 8840 15180 8840 0 _100_
rlabel metal2 7590 12852 7590 12852 0 _101_
rlabel metal4 9476 7072 9476 7072 0 _102_
rlabel metal2 15318 3468 15318 3468 0 _103_
rlabel metal1 16752 16422 16752 16422 0 _104_
rlabel metal1 17572 16694 17572 16694 0 _105_
rlabel metal1 8142 14382 8142 14382 0 _106_
rlabel metal1 9982 11220 9982 11220 0 _107_
rlabel metal1 10166 11254 10166 11254 0 _108_
rlabel metal2 5474 4284 5474 4284 0 _109_
rlabel metal3 3910 10268 3910 10268 0 _110_
rlabel metal2 5842 5134 5842 5134 0 _111_
rlabel metal2 9522 3196 9522 3196 0 _112_
rlabel metal1 2530 6222 2530 6222 0 _113_
rlabel metal2 18354 9129 18354 9129 0 _114_
rlabel metal1 4002 5712 4002 5712 0 _115_
rlabel metal1 15962 14382 15962 14382 0 _116_
rlabel metal1 15686 14518 15686 14518 0 _117_
rlabel metal1 7544 13430 7544 13430 0 _118_
rlabel metal2 10718 9248 10718 9248 0 _119_
rlabel metal1 17894 4250 17894 4250 0 _120_
rlabel metal1 8188 10506 8188 10506 0 _121_
rlabel metal1 1564 4114 1564 4114 0 _122_
rlabel metal1 14352 9622 14352 9622 0 _123_
rlabel metal1 14306 9452 14306 9452 0 _124_
rlabel metal1 12972 9554 12972 9554 0 _125_
rlabel metal2 13892 13396 13892 13396 0 _126_
rlabel metal1 5244 9078 5244 9078 0 _127_
rlabel metal1 9890 5134 9890 5134 0 _128_
rlabel metal1 4554 10166 4554 10166 0 _129_
rlabel via3 13915 15300 13915 15300 0 _130_
rlabel metal1 6532 13906 6532 13906 0 _131_
rlabel metal3 13662 8500 13662 8500 0 _132_
rlabel metal2 13662 6426 13662 6426 0 _133_
rlabel metal1 2208 10642 2208 10642 0 _134_
rlabel metal1 9154 2414 9154 2414 0 _135_
rlabel metal1 9200 15334 9200 15334 0 bloomFilter\[0\]
rlabel metal2 11730 12852 11730 12852 0 bloomFilter\[10\]
rlabel metal1 9338 12750 9338 12750 0 bloomFilter\[11\]
rlabel metal1 6532 8398 6532 8398 0 bloomFilter\[12\]
rlabel metal2 12190 15283 12190 15283 0 bloomFilter\[13\]
rlabel metal1 7280 8398 7280 8398 0 bloomFilter\[14\]
rlabel metal1 15870 13838 15870 13838 0 bloomFilter\[15\]
rlabel metal1 13754 14790 13754 14790 0 bloomFilter\[1\]
rlabel metal2 12466 7650 12466 7650 0 bloomFilter\[2\]
rlabel metal2 7130 11832 7130 11832 0 bloomFilter\[3\]
rlabel metal2 4416 9996 4416 9996 0 bloomFilter\[4\]
rlabel metal1 5060 4522 5060 4522 0 bloomFilter\[5\]
rlabel metal1 2254 12240 2254 12240 0 bloomFilter\[6\]
rlabel metal1 12328 9894 12328 9894 0 bloomFilter\[7\]
rlabel metal1 5888 5134 5888 5134 0 bloomFilter\[8\]
rlabel metal1 16652 12614 16652 12614 0 bloomFilter\[9\]
rlabel metal1 18262 2414 18262 2414 0 clk
rlabel via2 18446 6171 18446 6171 0 count[0]
rlabel metal2 8418 959 8418 959 0 count[10]
rlabel metal3 1142 15028 1142 15028 0 count[11]
rlabel metal3 820 6188 820 6188 0 count[12]
rlabel metal3 1142 18428 1142 18428 0 count[13]
rlabel metal1 18170 16762 18170 16762 0 count[14]
rlabel metal2 14214 1520 14214 1520 0 count[15]
rlabel metal3 820 2788 820 2788 0 count[1]
rlabel metal1 15640 17306 15640 17306 0 count[2]
rlabel metal1 18032 17306 18032 17306 0 count[3]
rlabel metal3 820 8908 820 8908 0 count[4]
rlabel metal2 4186 17595 4186 17595 0 count[5]
rlabel metal2 17434 1520 17434 1520 0 count[6]
rlabel metal2 46 1520 46 1520 0 count[7]
rlabel metal2 2622 959 2622 959 0 count[8]
rlabel metal1 6716 17306 6716 17306 0 count[9]
rlabel via2 18170 3451 18170 3451 0 enable
rlabel metal2 5842 1588 5842 1588 0 inputData[0]
rlabel metal3 18776 12308 18776 12308 0 inputData[1]
rlabel metal2 18262 15895 18262 15895 0 inputData[2]
rlabel metal1 9752 17170 9752 17170 0 inputData[3]
rlabel metal2 12282 18234 12282 18234 0 inputData[4]
rlabel metal2 11638 1588 11638 1588 0 inputData[5]
rlabel metal3 1142 12308 1142 12308 0 inputData[6]
rlabel metal1 2162 17204 2162 17204 0 inputData[7]
rlabel metal1 17066 5270 17066 5270 0 net1
rlabel metal1 1978 17000 1978 17000 0 net10
rlabel metal1 16606 8942 16606 8942 0 net11
rlabel metal1 18170 6290 18170 6290 0 net12
rlabel metal1 8556 2414 8556 2414 0 net13
rlabel via2 14122 12189 14122 12189 0 net14
rlabel metal2 1518 5916 1518 5916 0 net15
rlabel metal1 16744 16082 16744 16082 0 net16
rlabel via1 6578 12291 6578 12291 0 net17
rlabel metal1 12190 2482 12190 2482 0 net18
rlabel metal2 14030 12308 14030 12308 0 net19
rlabel metal2 14214 4794 14214 4794 0 net2
rlabel via2 2162 4165 2162 4165 0 net20
rlabel metal1 17250 17170 17250 17170 0 net21
rlabel metal1 3818 8466 3818 8466 0 net22
rlabel metal2 12650 15929 12650 15929 0 net23
rlabel metal1 15548 3094 15548 3094 0 net24
rlabel metal1 3864 2482 3864 2482 0 net25
rlabel metal1 4853 2346 4853 2346 0 net26
rlabel metal1 6946 12818 6946 12818 0 net27
rlabel metal1 2622 12682 2622 12682 0 net28
rlabel metal1 8602 9588 8602 9588 0 net29
rlabel metal1 15134 13328 15134 13328 0 net3
rlabel metal1 9154 2482 9154 2482 0 net30
rlabel metal1 15456 5338 15456 5338 0 net31
rlabel metal1 18216 12954 18216 12954 0 net4
rlabel metal2 2162 13073 2162 13073 0 net5
rlabel metal1 2116 4114 2116 4114 0 net6
rlabel metal2 15226 16558 15226 16558 0 net7
rlabel metal1 12788 2618 12788 2618 0 net8
rlabel metal2 5658 14518 5658 14518 0 net9
rlabel metal2 18170 9775 18170 9775 0 reset
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
